library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

ENTITY binaryToBCD is

	port( input: in std_logic_vector(15 downto 0);
			d1, d2, d3, d4: out std_logic_vector(3 downto 0)
	);
	
end ENTITY;

architecture behv of binaryToBCD is


	begin

		process(input)
		
			begin
			
			case input is
				    when "0000000000000000" => d1 <= "0000"; d2 <= "0000"; d3 <= "0000"; d4 <= "0000"; -- 0
    when "0000000000000001" => d1 <= "0001"; d2 <= "0000"; d3 <= "0000"; d4 <= "0000"; -- 1
    when "0000000000000010" => d1 <= "0010"; d2 <= "0000"; d3 <= "0000"; d4 <= "0000"; -- 2
    when "0000000000000011" => d1 <= "0011"; d2 <= "0000"; d3 <= "0000"; d4 <= "0000"; -- 3
    when "0000000000000100" => d1 <= "0100"; d2 <= "0000"; d3 <= "0000"; d4 <= "0000"; -- 4
    when "0000000000000101" => d1 <= "0101"; d2 <= "0000"; d3 <= "0000"; d4 <= "0000"; -- 5
    when "0000000000000110" => d1 <= "0110"; d2 <= "0000"; d3 <= "0000"; d4 <= "0000"; -- 6
    when "0000000000000111" => d1 <= "0111"; d2 <= "0000"; d3 <= "0000"; d4 <= "0000"; -- 7
    when "0000000000001000" => d1 <= "1000"; d2 <= "0000"; d3 <= "0000"; d4 <= "0000"; -- 8
    when "0000000000001001" => d1 <= "1001"; d2 <= "0000"; d3 <= "0000"; d4 <= "0000"; -- 9
    when "0000000000001010" => d1 <= "0000"; d2 <= "0001"; d3 <= "0000"; d4 <= "0000"; -- 10
    when "0000000000001011" => d1 <= "0001"; d2 <= "0001"; d3 <= "0000"; d4 <= "0000"; -- 11
    when "0000000000001100" => d1 <= "0010"; d2 <= "0001"; d3 <= "0000"; d4 <= "0000"; -- 12
    when "0000000000001101" => d1 <= "0011"; d2 <= "0001"; d3 <= "0000"; d4 <= "0000"; -- 13
    when "0000000000001110" => d1 <= "0100"; d2 <= "0001"; d3 <= "0000"; d4 <= "0000"; -- 14
    when "0000000000001111" => d1 <= "0101"; d2 <= "0001"; d3 <= "0000"; d4 <= "0000"; -- 15
    when "0000000000010000" => d1 <= "0110"; d2 <= "0001"; d3 <= "0000"; d4 <= "0000"; -- 16
    when "0000000000010001" => d1 <= "0111"; d2 <= "0001"; d3 <= "0000"; d4 <= "0000"; -- 17
    when "0000000000010010" => d1 <= "1000"; d2 <= "0001"; d3 <= "0000"; d4 <= "0000"; -- 18
    when "0000000000010011" => d1 <= "1001"; d2 <= "0001"; d3 <= "0000"; d4 <= "0000"; -- 19
    when "0000000000010100" => d1 <= "0000"; d2 <= "0010"; d3 <= "0000"; d4 <= "0000"; -- 20
    when "0000000000010101" => d1 <= "0001"; d2 <= "0010"; d3 <= "0000"; d4 <= "0000"; -- 21
    when "0000000000010110" => d1 <= "0010"; d2 <= "0010"; d3 <= "0000"; d4 <= "0000"; -- 22
    when "0000000000010111" => d1 <= "0011"; d2 <= "0010"; d3 <= "0000"; d4 <= "0000"; -- 23
    when "0000000000011000" => d1 <= "0100"; d2 <= "0010"; d3 <= "0000"; d4 <= "0000"; -- 24
    when "0000000000011001" => d1 <= "0101"; d2 <= "0010"; d3 <= "0000"; d4 <= "0000"; -- 25
    when "0000000000011010" => d1 <= "0110"; d2 <= "0010"; d3 <= "0000"; d4 <= "0000"; -- 26
    when "0000000000011011" => d1 <= "0111"; d2 <= "0010"; d3 <= "0000"; d4 <= "0000"; -- 27
    when "0000000000011100" => d1 <= "1000"; d2 <= "0010"; d3 <= "0000"; d4 <= "0000"; -- 28
    when "0000000000011101" => d1 <= "1001"; d2 <= "0010"; d3 <= "0000"; d4 <= "0000"; -- 29
    when "0000000000011110" => d1 <= "0000"; d2 <= "0011"; d3 <= "0000"; d4 <= "0000"; -- 30
    when "0000000000011111" => d1 <= "0001"; d2 <= "0011"; d3 <= "0000"; d4 <= "0000"; -- 31
    when "0000000000100000" => d1 <= "0010"; d2 <= "0011"; d3 <= "0000"; d4 <= "0000"; -- 32
    when "0000000000100001" => d1 <= "0011"; d2 <= "0011"; d3 <= "0000"; d4 <= "0000"; -- 33
    when "0000000000100010" => d1 <= "0100"; d2 <= "0011"; d3 <= "0000"; d4 <= "0000"; -- 34
    when "0000000000100011" => d1 <= "0101"; d2 <= "0011"; d3 <= "0000"; d4 <= "0000"; -- 35
    when "0000000000100100" => d1 <= "0110"; d2 <= "0011"; d3 <= "0000"; d4 <= "0000"; -- 36
    when "0000000000100101" => d1 <= "0111"; d2 <= "0011"; d3 <= "0000"; d4 <= "0000"; -- 37
    when "0000000000100110" => d1 <= "1000"; d2 <= "0011"; d3 <= "0000"; d4 <= "0000"; -- 38
    when "0000000000100111" => d1 <= "1001"; d2 <= "0011"; d3 <= "0000"; d4 <= "0000"; -- 39
    when "0000000000101000" => d1 <= "0000"; d2 <= "0100"; d3 <= "0000"; d4 <= "0000"; -- 40
    when "0000000000101001" => d1 <= "0001"; d2 <= "0100"; d3 <= "0000"; d4 <= "0000"; -- 41
    when "0000000000101010" => d1 <= "0010"; d2 <= "0100"; d3 <= "0000"; d4 <= "0000"; -- 42
    when "0000000000101011" => d1 <= "0011"; d2 <= "0100"; d3 <= "0000"; d4 <= "0000"; -- 43
    when "0000000000101100" => d1 <= "0100"; d2 <= "0100"; d3 <= "0000"; d4 <= "0000"; -- 44
    when "0000000000101101" => d1 <= "0101"; d2 <= "0100"; d3 <= "0000"; d4 <= "0000"; -- 45
    when "0000000000101110" => d1 <= "0110"; d2 <= "0100"; d3 <= "0000"; d4 <= "0000"; -- 46
    when "0000000000101111" => d1 <= "0111"; d2 <= "0100"; d3 <= "0000"; d4 <= "0000"; -- 47
    when "0000000000110000" => d1 <= "1000"; d2 <= "0100"; d3 <= "0000"; d4 <= "0000"; -- 48
    when "0000000000110001" => d1 <= "1001"; d2 <= "0100"; d3 <= "0000"; d4 <= "0000"; -- 49
    when "0000000000110010" => d1 <= "0000"; d2 <= "0101"; d3 <= "0000"; d4 <= "0000"; -- 50
    when "0000000000110011" => d1 <= "0001"; d2 <= "0101"; d3 <= "0000"; d4 <= "0000"; -- 51
    when "0000000000110100" => d1 <= "0010"; d2 <= "0101"; d3 <= "0000"; d4 <= "0000"; -- 52
    when "0000000000110101" => d1 <= "0011"; d2 <= "0101"; d3 <= "0000"; d4 <= "0000"; -- 53
    when "0000000000110110" => d1 <= "0100"; d2 <= "0101"; d3 <= "0000"; d4 <= "0000"; -- 54
    when "0000000000110111" => d1 <= "0101"; d2 <= "0101"; d3 <= "0000"; d4 <= "0000"; -- 55
    when "0000000000111000" => d1 <= "0110"; d2 <= "0101"; d3 <= "0000"; d4 <= "0000"; -- 56
    when "0000000000111001" => d1 <= "0111"; d2 <= "0101"; d3 <= "0000"; d4 <= "0000"; -- 57
    when "0000000000111010" => d1 <= "1000"; d2 <= "0101"; d3 <= "0000"; d4 <= "0000"; -- 58
    when "0000000000111011" => d1 <= "1001"; d2 <= "0101"; d3 <= "0000"; d4 <= "0000"; -- 59
    when "0000000000111100" => d1 <= "0000"; d2 <= "0110"; d3 <= "0000"; d4 <= "0000"; -- 60
    when "0000000000111101" => d1 <= "0001"; d2 <= "0110"; d3 <= "0000"; d4 <= "0000"; -- 61
    when "0000000000111110" => d1 <= "0010"; d2 <= "0110"; d3 <= "0000"; d4 <= "0000"; -- 62
    when "0000000000111111" => d1 <= "0011"; d2 <= "0110"; d3 <= "0000"; d4 <= "0000"; -- 63
    when "0000000001000000" => d1 <= "0100"; d2 <= "0110"; d3 <= "0000"; d4 <= "0000"; -- 64
    when "0000000001000001" => d1 <= "0101"; d2 <= "0110"; d3 <= "0000"; d4 <= "0000"; -- 65
    when "0000000001000010" => d1 <= "0110"; d2 <= "0110"; d3 <= "0000"; d4 <= "0000"; -- 66
    when "0000000001000011" => d1 <= "0111"; d2 <= "0110"; d3 <= "0000"; d4 <= "0000"; -- 67
    when "0000000001000100" => d1 <= "1000"; d2 <= "0110"; d3 <= "0000"; d4 <= "0000"; -- 68
    when "0000000001000101" => d1 <= "1001"; d2 <= "0110"; d3 <= "0000"; d4 <= "0000"; -- 69
    when "0000000001000110" => d1 <= "0000"; d2 <= "0111"; d3 <= "0000"; d4 <= "0000"; -- 70
    when "0000000001000111" => d1 <= "0001"; d2 <= "0111"; d3 <= "0000"; d4 <= "0000"; -- 71
    when "0000000001001000" => d1 <= "0010"; d2 <= "0111"; d3 <= "0000"; d4 <= "0000"; -- 72
    when "0000000001001001" => d1 <= "0011"; d2 <= "0111"; d3 <= "0000"; d4 <= "0000"; -- 73
    when "0000000001001010" => d1 <= "0100"; d2 <= "0111"; d3 <= "0000"; d4 <= "0000"; -- 74
    when "0000000001001011" => d1 <= "0101"; d2 <= "0111"; d3 <= "0000"; d4 <= "0000"; -- 75
    when "0000000001001100" => d1 <= "0110"; d2 <= "0111"; d3 <= "0000"; d4 <= "0000"; -- 76
    when "0000000001001101" => d1 <= "0111"; d2 <= "0111"; d3 <= "0000"; d4 <= "0000"; -- 77
    when "0000000001001110" => d1 <= "1000"; d2 <= "0111"; d3 <= "0000"; d4 <= "0000"; -- 78
    when "0000000001001111" => d1 <= "1001"; d2 <= "0111"; d3 <= "0000"; d4 <= "0000"; -- 79
    when "0000000001010000" => d1 <= "0000"; d2 <= "1000"; d3 <= "0000"; d4 <= "0000"; -- 80
    when "0000000001010001" => d1 <= "0001"; d2 <= "1000"; d3 <= "0000"; d4 <= "0000"; -- 81
    when "0000000001010010" => d1 <= "0010"; d2 <= "1000"; d3 <= "0000"; d4 <= "0000"; -- 82
    when "0000000001010011" => d1 <= "0011"; d2 <= "1000"; d3 <= "0000"; d4 <= "0000"; -- 83
    when "0000000001010100" => d1 <= "0100"; d2 <= "1000"; d3 <= "0000"; d4 <= "0000"; -- 84
    when "0000000001010101" => d1 <= "0101"; d2 <= "1000"; d3 <= "0000"; d4 <= "0000"; -- 85
    when "0000000001010110" => d1 <= "0110"; d2 <= "1000"; d3 <= "0000"; d4 <= "0000"; -- 86
    when "0000000001010111" => d1 <= "0111"; d2 <= "1000"; d3 <= "0000"; d4 <= "0000"; -- 87
    when "0000000001011000" => d1 <= "1000"; d2 <= "1000"; d3 <= "0000"; d4 <= "0000"; -- 88
    when "0000000001011001" => d1 <= "1001"; d2 <= "1000"; d3 <= "0000"; d4 <= "0000"; -- 89
    when "0000000001011010" => d1 <= "0000"; d2 <= "1001"; d3 <= "0000"; d4 <= "0000"; -- 90
    when "0000000001011011" => d1 <= "0001"; d2 <= "1001"; d3 <= "0000"; d4 <= "0000"; -- 91
    when "0000000001011100" => d1 <= "0010"; d2 <= "1001"; d3 <= "0000"; d4 <= "0000"; -- 92
    when "0000000001011101" => d1 <= "0011"; d2 <= "1001"; d3 <= "0000"; d4 <= "0000"; -- 93
    when "0000000001011110" => d1 <= "0100"; d2 <= "1001"; d3 <= "0000"; d4 <= "0000"; -- 94
    when "0000000001011111" => d1 <= "0101"; d2 <= "1001"; d3 <= "0000"; d4 <= "0000"; -- 95
    when "0000000001100000" => d1 <= "0110"; d2 <= "1001"; d3 <= "0000"; d4 <= "0000"; -- 96
    when "0000000001100001" => d1 <= "0111"; d2 <= "1001"; d3 <= "0000"; d4 <= "0000"; -- 97
    when "0000000001100010" => d1 <= "1000"; d2 <= "1001"; d3 <= "0000"; d4 <= "0000"; -- 98
    when "0000000001100011" => d1 <= "1001"; d2 <= "1001"; d3 <= "0000"; d4 <= "0000"; -- 99
    when "0000000001100100" => d1 <= "0000"; d2 <= "0000"; d3 <= "0001"; d4 <= "0000"; -- 100
    when "0000000001100101" => d1 <= "0001"; d2 <= "0000"; d3 <= "0001"; d4 <= "0000"; -- 101
    when "0000000001100110" => d1 <= "0010"; d2 <= "0000"; d3 <= "0001"; d4 <= "0000"; -- 102
    when "0000000001100111" => d1 <= "0011"; d2 <= "0000"; d3 <= "0001"; d4 <= "0000"; -- 103
    when "0000000001101000" => d1 <= "0100"; d2 <= "0000"; d3 <= "0001"; d4 <= "0000"; -- 104
    when "0000000001101001" => d1 <= "0101"; d2 <= "0000"; d3 <= "0001"; d4 <= "0000"; -- 105
    when "0000000001101010" => d1 <= "0110"; d2 <= "0000"; d3 <= "0001"; d4 <= "0000"; -- 106
    when "0000000001101011" => d1 <= "0111"; d2 <= "0000"; d3 <= "0001"; d4 <= "0000"; -- 107
    when "0000000001101100" => d1 <= "1000"; d2 <= "0000"; d3 <= "0001"; d4 <= "0000"; -- 108
    when "0000000001101101" => d1 <= "1001"; d2 <= "0000"; d3 <= "0001"; d4 <= "0000"; -- 109
    when "0000000001101110" => d1 <= "0000"; d2 <= "0001"; d3 <= "0001"; d4 <= "0000"; -- 110
    when "0000000001101111" => d1 <= "0001"; d2 <= "0001"; d3 <= "0001"; d4 <= "0000"; -- 111
    when "0000000001110000" => d1 <= "0010"; d2 <= "0001"; d3 <= "0001"; d4 <= "0000"; -- 112
    when "0000000001110001" => d1 <= "0011"; d2 <= "0001"; d3 <= "0001"; d4 <= "0000"; -- 113
    when "0000000001110010" => d1 <= "0100"; d2 <= "0001"; d3 <= "0001"; d4 <= "0000"; -- 114
    when "0000000001110011" => d1 <= "0101"; d2 <= "0001"; d3 <= "0001"; d4 <= "0000"; -- 115
    when "0000000001110100" => d1 <= "0110"; d2 <= "0001"; d3 <= "0001"; d4 <= "0000"; -- 116
    when "0000000001110101" => d1 <= "0111"; d2 <= "0001"; d3 <= "0001"; d4 <= "0000"; -- 117
    when "0000000001110110" => d1 <= "1000"; d2 <= "0001"; d3 <= "0001"; d4 <= "0000"; -- 118
    when "0000000001110111" => d1 <= "1001"; d2 <= "0001"; d3 <= "0001"; d4 <= "0000"; -- 119
    when "0000000001111000" => d1 <= "0000"; d2 <= "0010"; d3 <= "0001"; d4 <= "0000"; -- 120
    when "0000000001111001" => d1 <= "0001"; d2 <= "0010"; d3 <= "0001"; d4 <= "0000"; -- 121
    when "0000000001111010" => d1 <= "0010"; d2 <= "0010"; d3 <= "0001"; d4 <= "0000"; -- 122
    when "0000000001111011" => d1 <= "0011"; d2 <= "0010"; d3 <= "0001"; d4 <= "0000"; -- 123
    when "0000000001111100" => d1 <= "0100"; d2 <= "0010"; d3 <= "0001"; d4 <= "0000"; -- 124
    when "0000000001111101" => d1 <= "0101"; d2 <= "0010"; d3 <= "0001"; d4 <= "0000"; -- 125
    when "0000000001111110" => d1 <= "0110"; d2 <= "0010"; d3 <= "0001"; d4 <= "0000"; -- 126
    when "0000000001111111" => d1 <= "0111"; d2 <= "0010"; d3 <= "0001"; d4 <= "0000"; -- 127
    when "0000000010000000" => d1 <= "1000"; d2 <= "0010"; d3 <= "0001"; d4 <= "0000"; -- 128
    when "0000000010000001" => d1 <= "1001"; d2 <= "0010"; d3 <= "0001"; d4 <= "0000"; -- 129
    when "0000000010000010" => d1 <= "0000"; d2 <= "0011"; d3 <= "0001"; d4 <= "0000"; -- 130
    when "0000000010000011" => d1 <= "0001"; d2 <= "0011"; d3 <= "0001"; d4 <= "0000"; -- 131
    when "0000000010000100" => d1 <= "0010"; d2 <= "0011"; d3 <= "0001"; d4 <= "0000"; -- 132
    when "0000000010000101" => d1 <= "0011"; d2 <= "0011"; d3 <= "0001"; d4 <= "0000"; -- 133
    when "0000000010000110" => d1 <= "0100"; d2 <= "0011"; d3 <= "0001"; d4 <= "0000"; -- 134
    when "0000000010000111" => d1 <= "0101"; d2 <= "0011"; d3 <= "0001"; d4 <= "0000"; -- 135
    when "0000000010001000" => d1 <= "0110"; d2 <= "0011"; d3 <= "0001"; d4 <= "0000"; -- 136
    when "0000000010001001" => d1 <= "0111"; d2 <= "0011"; d3 <= "0001"; d4 <= "0000"; -- 137
    when "0000000010001010" => d1 <= "1000"; d2 <= "0011"; d3 <= "0001"; d4 <= "0000"; -- 138
    when "0000000010001011" => d1 <= "1001"; d2 <= "0011"; d3 <= "0001"; d4 <= "0000"; -- 139
    when "0000000010001100" => d1 <= "0000"; d2 <= "0100"; d3 <= "0001"; d4 <= "0000"; -- 140
    when "0000000010001101" => d1 <= "0001"; d2 <= "0100"; d3 <= "0001"; d4 <= "0000"; -- 141
    when "0000000010001110" => d1 <= "0010"; d2 <= "0100"; d3 <= "0001"; d4 <= "0000"; -- 142
    when "0000000010001111" => d1 <= "0011"; d2 <= "0100"; d3 <= "0001"; d4 <= "0000"; -- 143
    when "0000000010010000" => d1 <= "0100"; d2 <= "0100"; d3 <= "0001"; d4 <= "0000"; -- 144
    when "0000000010010001" => d1 <= "0101"; d2 <= "0100"; d3 <= "0001"; d4 <= "0000"; -- 145
    when "0000000010010010" => d1 <= "0110"; d2 <= "0100"; d3 <= "0001"; d4 <= "0000"; -- 146
    when "0000000010010011" => d1 <= "0111"; d2 <= "0100"; d3 <= "0001"; d4 <= "0000"; -- 147
    when "0000000010010100" => d1 <= "1000"; d2 <= "0100"; d3 <= "0001"; d4 <= "0000"; -- 148
    when "0000000010010101" => d1 <= "1001"; d2 <= "0100"; d3 <= "0001"; d4 <= "0000"; -- 149
    when "0000000010010110" => d1 <= "0000"; d2 <= "0101"; d3 <= "0001"; d4 <= "0000"; -- 150
    when "0000000010010111" => d1 <= "0001"; d2 <= "0101"; d3 <= "0001"; d4 <= "0000"; -- 151
    when "0000000010011000" => d1 <= "0010"; d2 <= "0101"; d3 <= "0001"; d4 <= "0000"; -- 152
    when "0000000010011001" => d1 <= "0011"; d2 <= "0101"; d3 <= "0001"; d4 <= "0000"; -- 153
    when "0000000010011010" => d1 <= "0100"; d2 <= "0101"; d3 <= "0001"; d4 <= "0000"; -- 154
    when "0000000010011011" => d1 <= "0101"; d2 <= "0101"; d3 <= "0001"; d4 <= "0000"; -- 155
    when "0000000010011100" => d1 <= "0110"; d2 <= "0101"; d3 <= "0001"; d4 <= "0000"; -- 156
    when "0000000010011101" => d1 <= "0111"; d2 <= "0101"; d3 <= "0001"; d4 <= "0000"; -- 157
    when "0000000010011110" => d1 <= "1000"; d2 <= "0101"; d3 <= "0001"; d4 <= "0000"; -- 158
    when "0000000010011111" => d1 <= "1001"; d2 <= "0101"; d3 <= "0001"; d4 <= "0000"; -- 159
    when "0000000010100000" => d1 <= "0000"; d2 <= "0110"; d3 <= "0001"; d4 <= "0000"; -- 160
    when "0000000010100001" => d1 <= "0001"; d2 <= "0110"; d3 <= "0001"; d4 <= "0000"; -- 161
    when "0000000010100010" => d1 <= "0010"; d2 <= "0110"; d3 <= "0001"; d4 <= "0000"; -- 162
    when "0000000010100011" => d1 <= "0011"; d2 <= "0110"; d3 <= "0001"; d4 <= "0000"; -- 163
    when "0000000010100100" => d1 <= "0100"; d2 <= "0110"; d3 <= "0001"; d4 <= "0000"; -- 164
    when "0000000010100101" => d1 <= "0101"; d2 <= "0110"; d3 <= "0001"; d4 <= "0000"; -- 165
    when "0000000010100110" => d1 <= "0110"; d2 <= "0110"; d3 <= "0001"; d4 <= "0000"; -- 166
    when "0000000010100111" => d1 <= "0111"; d2 <= "0110"; d3 <= "0001"; d4 <= "0000"; -- 167
    when "0000000010101000" => d1 <= "1000"; d2 <= "0110"; d3 <= "0001"; d4 <= "0000"; -- 168
    when "0000000010101001" => d1 <= "1001"; d2 <= "0110"; d3 <= "0001"; d4 <= "0000"; -- 169
    when "0000000010101010" => d1 <= "0000"; d2 <= "0111"; d3 <= "0001"; d4 <= "0000"; -- 170
    when "0000000010101011" => d1 <= "0001"; d2 <= "0111"; d3 <= "0001"; d4 <= "0000"; -- 171
    when "0000000010101100" => d1 <= "0010"; d2 <= "0111"; d3 <= "0001"; d4 <= "0000"; -- 172
    when "0000000010101101" => d1 <= "0011"; d2 <= "0111"; d3 <= "0001"; d4 <= "0000"; -- 173
    when "0000000010101110" => d1 <= "0100"; d2 <= "0111"; d3 <= "0001"; d4 <= "0000"; -- 174
    when "0000000010101111" => d1 <= "0101"; d2 <= "0111"; d3 <= "0001"; d4 <= "0000"; -- 175
    when "0000000010110000" => d1 <= "0110"; d2 <= "0111"; d3 <= "0001"; d4 <= "0000"; -- 176
    when "0000000010110001" => d1 <= "0111"; d2 <= "0111"; d3 <= "0001"; d4 <= "0000"; -- 177
    when "0000000010110010" => d1 <= "1000"; d2 <= "0111"; d3 <= "0001"; d4 <= "0000"; -- 178
    when "0000000010110011" => d1 <= "1001"; d2 <= "0111"; d3 <= "0001"; d4 <= "0000"; -- 179
    when "0000000010110100" => d1 <= "0000"; d2 <= "1000"; d3 <= "0001"; d4 <= "0000"; -- 180
    when "0000000010110101" => d1 <= "0001"; d2 <= "1000"; d3 <= "0001"; d4 <= "0000"; -- 181
    when "0000000010110110" => d1 <= "0010"; d2 <= "1000"; d3 <= "0001"; d4 <= "0000"; -- 182
    when "0000000010110111" => d1 <= "0011"; d2 <= "1000"; d3 <= "0001"; d4 <= "0000"; -- 183
    when "0000000010111000" => d1 <= "0100"; d2 <= "1000"; d3 <= "0001"; d4 <= "0000"; -- 184
    when "0000000010111001" => d1 <= "0101"; d2 <= "1000"; d3 <= "0001"; d4 <= "0000"; -- 185
    when "0000000010111010" => d1 <= "0110"; d2 <= "1000"; d3 <= "0001"; d4 <= "0000"; -- 186
    when "0000000010111011" => d1 <= "0111"; d2 <= "1000"; d3 <= "0001"; d4 <= "0000"; -- 187
    when "0000000010111100" => d1 <= "1000"; d2 <= "1000"; d3 <= "0001"; d4 <= "0000"; -- 188
    when "0000000010111101" => d1 <= "1001"; d2 <= "1000"; d3 <= "0001"; d4 <= "0000"; -- 189
    when "0000000010111110" => d1 <= "0000"; d2 <= "1001"; d3 <= "0001"; d4 <= "0000"; -- 190
    when "0000000010111111" => d1 <= "0001"; d2 <= "1001"; d3 <= "0001"; d4 <= "0000"; -- 191
    when "0000000011000000" => d1 <= "0010"; d2 <= "1001"; d3 <= "0001"; d4 <= "0000"; -- 192
    when "0000000011000001" => d1 <= "0011"; d2 <= "1001"; d3 <= "0001"; d4 <= "0000"; -- 193
    when "0000000011000010" => d1 <= "0100"; d2 <= "1001"; d3 <= "0001"; d4 <= "0000"; -- 194
    when "0000000011000011" => d1 <= "0101"; d2 <= "1001"; d3 <= "0001"; d4 <= "0000"; -- 195
    when "0000000011000100" => d1 <= "0110"; d2 <= "1001"; d3 <= "0001"; d4 <= "0000"; -- 196
    when "0000000011000101" => d1 <= "0111"; d2 <= "1001"; d3 <= "0001"; d4 <= "0000"; -- 197
    when "0000000011000110" => d1 <= "1000"; d2 <= "1001"; d3 <= "0001"; d4 <= "0000"; -- 198
    when "0000000011000111" => d1 <= "1001"; d2 <= "1001"; d3 <= "0001"; d4 <= "0000"; -- 199
    when "0000000011001000" => d1 <= "0000"; d2 <= "0000"; d3 <= "0010"; d4 <= "0000"; -- 200
    when "0000000011001001" => d1 <= "0001"; d2 <= "0000"; d3 <= "0010"; d4 <= "0000"; -- 201
    when "0000000011001010" => d1 <= "0010"; d2 <= "0000"; d3 <= "0010"; d4 <= "0000"; -- 202
    when "0000000011001011" => d1 <= "0011"; d2 <= "0000"; d3 <= "0010"; d4 <= "0000"; -- 203
    when "0000000011001100" => d1 <= "0100"; d2 <= "0000"; d3 <= "0010"; d4 <= "0000"; -- 204
    when "0000000011001101" => d1 <= "0101"; d2 <= "0000"; d3 <= "0010"; d4 <= "0000"; -- 205
    when "0000000011001110" => d1 <= "0110"; d2 <= "0000"; d3 <= "0010"; d4 <= "0000"; -- 206
    when "0000000011001111" => d1 <= "0111"; d2 <= "0000"; d3 <= "0010"; d4 <= "0000"; -- 207
    when "0000000011010000" => d1 <= "1000"; d2 <= "0000"; d3 <= "0010"; d4 <= "0000"; -- 208
    when "0000000011010001" => d1 <= "1001"; d2 <= "0000"; d3 <= "0010"; d4 <= "0000"; -- 209
    when "0000000011010010" => d1 <= "0000"; d2 <= "0001"; d3 <= "0010"; d4 <= "0000"; -- 210
    when "0000000011010011" => d1 <= "0001"; d2 <= "0001"; d3 <= "0010"; d4 <= "0000"; -- 211
    when "0000000011010100" => d1 <= "0010"; d2 <= "0001"; d3 <= "0010"; d4 <= "0000"; -- 212
    when "0000000011010101" => d1 <= "0011"; d2 <= "0001"; d3 <= "0010"; d4 <= "0000"; -- 213
    when "0000000011010110" => d1 <= "0100"; d2 <= "0001"; d3 <= "0010"; d4 <= "0000"; -- 214
    when "0000000011010111" => d1 <= "0101"; d2 <= "0001"; d3 <= "0010"; d4 <= "0000"; -- 215
    when "0000000011011000" => d1 <= "0110"; d2 <= "0001"; d3 <= "0010"; d4 <= "0000"; -- 216
    when "0000000011011001" => d1 <= "0111"; d2 <= "0001"; d3 <= "0010"; d4 <= "0000"; -- 217
    when "0000000011011010" => d1 <= "1000"; d2 <= "0001"; d3 <= "0010"; d4 <= "0000"; -- 218
    when "0000000011011011" => d1 <= "1001"; d2 <= "0001"; d3 <= "0010"; d4 <= "0000"; -- 219
    when "0000000011011100" => d1 <= "0000"; d2 <= "0010"; d3 <= "0010"; d4 <= "0000"; -- 220
    when "0000000011011101" => d1 <= "0001"; d2 <= "0010"; d3 <= "0010"; d4 <= "0000"; -- 221
    when "0000000011011110" => d1 <= "0010"; d2 <= "0010"; d3 <= "0010"; d4 <= "0000"; -- 222
    when "0000000011011111" => d1 <= "0011"; d2 <= "0010"; d3 <= "0010"; d4 <= "0000"; -- 223
    when "0000000011100000" => d1 <= "0100"; d2 <= "0010"; d3 <= "0010"; d4 <= "0000"; -- 224
    when "0000000011100001" => d1 <= "0101"; d2 <= "0010"; d3 <= "0010"; d4 <= "0000"; -- 225
    when "0000000011100010" => d1 <= "0110"; d2 <= "0010"; d3 <= "0010"; d4 <= "0000"; -- 226
    when "0000000011100011" => d1 <= "0111"; d2 <= "0010"; d3 <= "0010"; d4 <= "0000"; -- 227
    when "0000000011100100" => d1 <= "1000"; d2 <= "0010"; d3 <= "0010"; d4 <= "0000"; -- 228
    when "0000000011100101" => d1 <= "1001"; d2 <= "0010"; d3 <= "0010"; d4 <= "0000"; -- 229
    when "0000000011100110" => d1 <= "0000"; d2 <= "0011"; d3 <= "0010"; d4 <= "0000"; -- 230
    when "0000000011100111" => d1 <= "0001"; d2 <= "0011"; d3 <= "0010"; d4 <= "0000"; -- 231
    when "0000000011101000" => d1 <= "0010"; d2 <= "0011"; d3 <= "0010"; d4 <= "0000"; -- 232
    when "0000000011101001" => d1 <= "0011"; d2 <= "0011"; d3 <= "0010"; d4 <= "0000"; -- 233
    when "0000000011101010" => d1 <= "0100"; d2 <= "0011"; d3 <= "0010"; d4 <= "0000"; -- 234
    when "0000000011101011" => d1 <= "0101"; d2 <= "0011"; d3 <= "0010"; d4 <= "0000"; -- 235
    when "0000000011101100" => d1 <= "0110"; d2 <= "0011"; d3 <= "0010"; d4 <= "0000"; -- 236
    when "0000000011101101" => d1 <= "0111"; d2 <= "0011"; d3 <= "0010"; d4 <= "0000"; -- 237
    when "0000000011101110" => d1 <= "1000"; d2 <= "0011"; d3 <= "0010"; d4 <= "0000"; -- 238
    when "0000000011101111" => d1 <= "1001"; d2 <= "0011"; d3 <= "0010"; d4 <= "0000"; -- 239
    when "0000000011110000" => d1 <= "0000"; d2 <= "0100"; d3 <= "0010"; d4 <= "0000"; -- 240
    when "0000000011110001" => d1 <= "0001"; d2 <= "0100"; d3 <= "0010"; d4 <= "0000"; -- 241
    when "0000000011110010" => d1 <= "0010"; d2 <= "0100"; d3 <= "0010"; d4 <= "0000"; -- 242
    when "0000000011110011" => d1 <= "0011"; d2 <= "0100"; d3 <= "0010"; d4 <= "0000"; -- 243
    when "0000000011110100" => d1 <= "0100"; d2 <= "0100"; d3 <= "0010"; d4 <= "0000"; -- 244
    when "0000000011110101" => d1 <= "0101"; d2 <= "0100"; d3 <= "0010"; d4 <= "0000"; -- 245
    when "0000000011110110" => d1 <= "0110"; d2 <= "0100"; d3 <= "0010"; d4 <= "0000"; -- 246
    when "0000000011110111" => d1 <= "0111"; d2 <= "0100"; d3 <= "0010"; d4 <= "0000"; -- 247
    when "0000000011111000" => d1 <= "1000"; d2 <= "0100"; d3 <= "0010"; d4 <= "0000"; -- 248
    when "0000000011111001" => d1 <= "1001"; d2 <= "0100"; d3 <= "0010"; d4 <= "0000"; -- 249
    when "0000000011111010" => d1 <= "0000"; d2 <= "0101"; d3 <= "0010"; d4 <= "0000"; -- 250
    when "0000000011111011" => d1 <= "0001"; d2 <= "0101"; d3 <= "0010"; d4 <= "0000"; -- 251
    when "0000000011111100" => d1 <= "0010"; d2 <= "0101"; d3 <= "0010"; d4 <= "0000"; -- 252
    when "0000000011111101" => d1 <= "0011"; d2 <= "0101"; d3 <= "0010"; d4 <= "0000"; -- 253
    when "0000000011111110" => d1 <= "0100"; d2 <= "0101"; d3 <= "0010"; d4 <= "0000"; -- 254
    when "0000000011111111" => d1 <= "0101"; d2 <= "0101"; d3 <= "0010"; d4 <= "0000"; -- 255
    when "0000000100000000" => d1 <= "0110"; d2 <= "0101"; d3 <= "0010"; d4 <= "0000"; -- 256
    when "0000000100000001" => d1 <= "0111"; d2 <= "0101"; d3 <= "0010"; d4 <= "0000"; -- 257
    when "0000000100000010" => d1 <= "1000"; d2 <= "0101"; d3 <= "0010"; d4 <= "0000"; -- 258
    when "0000000100000011" => d1 <= "1001"; d2 <= "0101"; d3 <= "0010"; d4 <= "0000"; -- 259
    when "0000000100000100" => d1 <= "0000"; d2 <= "0110"; d3 <= "0010"; d4 <= "0000"; -- 260
    when "0000000100000101" => d1 <= "0001"; d2 <= "0110"; d3 <= "0010"; d4 <= "0000"; -- 261
    when "0000000100000110" => d1 <= "0010"; d2 <= "0110"; d3 <= "0010"; d4 <= "0000"; -- 262
    when "0000000100000111" => d1 <= "0011"; d2 <= "0110"; d3 <= "0010"; d4 <= "0000"; -- 263
    when "0000000100001000" => d1 <= "0100"; d2 <= "0110"; d3 <= "0010"; d4 <= "0000"; -- 264
    when "0000000100001001" => d1 <= "0101"; d2 <= "0110"; d3 <= "0010"; d4 <= "0000"; -- 265
    when "0000000100001010" => d1 <= "0110"; d2 <= "0110"; d3 <= "0010"; d4 <= "0000"; -- 266
    when "0000000100001011" => d1 <= "0111"; d2 <= "0110"; d3 <= "0010"; d4 <= "0000"; -- 267
    when "0000000100001100" => d1 <= "1000"; d2 <= "0110"; d3 <= "0010"; d4 <= "0000"; -- 268
    when "0000000100001101" => d1 <= "1001"; d2 <= "0110"; d3 <= "0010"; d4 <= "0000"; -- 269
    when "0000000100001110" => d1 <= "0000"; d2 <= "0111"; d3 <= "0010"; d4 <= "0000"; -- 270
    when "0000000100001111" => d1 <= "0001"; d2 <= "0111"; d3 <= "0010"; d4 <= "0000"; -- 271
    when "0000000100010000" => d1 <= "0010"; d2 <= "0111"; d3 <= "0010"; d4 <= "0000"; -- 272
    when "0000000100010001" => d1 <= "0011"; d2 <= "0111"; d3 <= "0010"; d4 <= "0000"; -- 273
    when "0000000100010010" => d1 <= "0100"; d2 <= "0111"; d3 <= "0010"; d4 <= "0000"; -- 274
    when "0000000100010011" => d1 <= "0101"; d2 <= "0111"; d3 <= "0010"; d4 <= "0000"; -- 275
    when "0000000100010100" => d1 <= "0110"; d2 <= "0111"; d3 <= "0010"; d4 <= "0000"; -- 276
    when "0000000100010101" => d1 <= "0111"; d2 <= "0111"; d3 <= "0010"; d4 <= "0000"; -- 277
    when "0000000100010110" => d1 <= "1000"; d2 <= "0111"; d3 <= "0010"; d4 <= "0000"; -- 278
    when "0000000100010111" => d1 <= "1001"; d2 <= "0111"; d3 <= "0010"; d4 <= "0000"; -- 279
    when "0000000100011000" => d1 <= "0000"; d2 <= "1000"; d3 <= "0010"; d4 <= "0000"; -- 280
    when "0000000100011001" => d1 <= "0001"; d2 <= "1000"; d3 <= "0010"; d4 <= "0000"; -- 281
    when "0000000100011010" => d1 <= "0010"; d2 <= "1000"; d3 <= "0010"; d4 <= "0000"; -- 282
    when "0000000100011011" => d1 <= "0011"; d2 <= "1000"; d3 <= "0010"; d4 <= "0000"; -- 283
    when "0000000100011100" => d1 <= "0100"; d2 <= "1000"; d3 <= "0010"; d4 <= "0000"; -- 284
    when "0000000100011101" => d1 <= "0101"; d2 <= "1000"; d3 <= "0010"; d4 <= "0000"; -- 285
    when "0000000100011110" => d1 <= "0110"; d2 <= "1000"; d3 <= "0010"; d4 <= "0000"; -- 286
    when "0000000100011111" => d1 <= "0111"; d2 <= "1000"; d3 <= "0010"; d4 <= "0000"; -- 287
    when "0000000100100000" => d1 <= "1000"; d2 <= "1000"; d3 <= "0010"; d4 <= "0000"; -- 288
    when "0000000100100001" => d1 <= "1001"; d2 <= "1000"; d3 <= "0010"; d4 <= "0000"; -- 289
    when "0000000100100010" => d1 <= "0000"; d2 <= "1001"; d3 <= "0010"; d4 <= "0000"; -- 290
    when "0000000100100011" => d1 <= "0001"; d2 <= "1001"; d3 <= "0010"; d4 <= "0000"; -- 291
    when "0000000100100100" => d1 <= "0010"; d2 <= "1001"; d3 <= "0010"; d4 <= "0000"; -- 292
    when "0000000100100101" => d1 <= "0011"; d2 <= "1001"; d3 <= "0010"; d4 <= "0000"; -- 293
    when "0000000100100110" => d1 <= "0100"; d2 <= "1001"; d3 <= "0010"; d4 <= "0000"; -- 294
    when "0000000100100111" => d1 <= "0101"; d2 <= "1001"; d3 <= "0010"; d4 <= "0000"; -- 295
    when "0000000100101000" => d1 <= "0110"; d2 <= "1001"; d3 <= "0010"; d4 <= "0000"; -- 296
    when "0000000100101001" => d1 <= "0111"; d2 <= "1001"; d3 <= "0010"; d4 <= "0000"; -- 297
    when "0000000100101010" => d1 <= "1000"; d2 <= "1001"; d3 <= "0010"; d4 <= "0000"; -- 298
    when "0000000100101011" => d1 <= "1001"; d2 <= "1001"; d3 <= "0010"; d4 <= "0000"; -- 299
    when "0000000100101100" => d1 <= "0000"; d2 <= "0000"; d3 <= "0011"; d4 <= "0000"; -- 300
    when "0000000100101101" => d1 <= "0001"; d2 <= "0000"; d3 <= "0011"; d4 <= "0000"; -- 301
    when "0000000100101110" => d1 <= "0010"; d2 <= "0000"; d3 <= "0011"; d4 <= "0000"; -- 302
    when "0000000100101111" => d1 <= "0011"; d2 <= "0000"; d3 <= "0011"; d4 <= "0000"; -- 303
    when "0000000100110000" => d1 <= "0100"; d2 <= "0000"; d3 <= "0011"; d4 <= "0000"; -- 304
    when "0000000100110001" => d1 <= "0101"; d2 <= "0000"; d3 <= "0011"; d4 <= "0000"; -- 305
    when "0000000100110010" => d1 <= "0110"; d2 <= "0000"; d3 <= "0011"; d4 <= "0000"; -- 306
    when "0000000100110011" => d1 <= "0111"; d2 <= "0000"; d3 <= "0011"; d4 <= "0000"; -- 307
    when "0000000100110100" => d1 <= "1000"; d2 <= "0000"; d3 <= "0011"; d4 <= "0000"; -- 308
    when "0000000100110101" => d1 <= "1001"; d2 <= "0000"; d3 <= "0011"; d4 <= "0000"; -- 309
    when "0000000100110110" => d1 <= "0000"; d2 <= "0001"; d3 <= "0011"; d4 <= "0000"; -- 310
    when "0000000100110111" => d1 <= "0001"; d2 <= "0001"; d3 <= "0011"; d4 <= "0000"; -- 311
    when "0000000100111000" => d1 <= "0010"; d2 <= "0001"; d3 <= "0011"; d4 <= "0000"; -- 312
    when "0000000100111001" => d1 <= "0011"; d2 <= "0001"; d3 <= "0011"; d4 <= "0000"; -- 313
    when "0000000100111010" => d1 <= "0100"; d2 <= "0001"; d3 <= "0011"; d4 <= "0000"; -- 314
    when "0000000100111011" => d1 <= "0101"; d2 <= "0001"; d3 <= "0011"; d4 <= "0000"; -- 315
    when "0000000100111100" => d1 <= "0110"; d2 <= "0001"; d3 <= "0011"; d4 <= "0000"; -- 316
    when "0000000100111101" => d1 <= "0111"; d2 <= "0001"; d3 <= "0011"; d4 <= "0000"; -- 317
    when "0000000100111110" => d1 <= "1000"; d2 <= "0001"; d3 <= "0011"; d4 <= "0000"; -- 318
    when "0000000100111111" => d1 <= "1001"; d2 <= "0001"; d3 <= "0011"; d4 <= "0000"; -- 319
    when "0000000101000000" => d1 <= "0000"; d2 <= "0010"; d3 <= "0011"; d4 <= "0000"; -- 320
    when "0000000101000001" => d1 <= "0001"; d2 <= "0010"; d3 <= "0011"; d4 <= "0000"; -- 321
    when "0000000101000010" => d1 <= "0010"; d2 <= "0010"; d3 <= "0011"; d4 <= "0000"; -- 322
    when "0000000101000011" => d1 <= "0011"; d2 <= "0010"; d3 <= "0011"; d4 <= "0000"; -- 323
    when "0000000101000100" => d1 <= "0100"; d2 <= "0010"; d3 <= "0011"; d4 <= "0000"; -- 324
    when "0000000101000101" => d1 <= "0101"; d2 <= "0010"; d3 <= "0011"; d4 <= "0000"; -- 325
    when "0000000101000110" => d1 <= "0110"; d2 <= "0010"; d3 <= "0011"; d4 <= "0000"; -- 326
    when "0000000101000111" => d1 <= "0111"; d2 <= "0010"; d3 <= "0011"; d4 <= "0000"; -- 327
    when "0000000101001000" => d1 <= "1000"; d2 <= "0010"; d3 <= "0011"; d4 <= "0000"; -- 328
    when "0000000101001001" => d1 <= "1001"; d2 <= "0010"; d3 <= "0011"; d4 <= "0000"; -- 329
    when "0000000101001010" => d1 <= "0000"; d2 <= "0011"; d3 <= "0011"; d4 <= "0000"; -- 330
    when "0000000101001011" => d1 <= "0001"; d2 <= "0011"; d3 <= "0011"; d4 <= "0000"; -- 331
    when "0000000101001100" => d1 <= "0010"; d2 <= "0011"; d3 <= "0011"; d4 <= "0000"; -- 332
    when "0000000101001101" => d1 <= "0011"; d2 <= "0011"; d3 <= "0011"; d4 <= "0000"; -- 333
    when "0000000101001110" => d1 <= "0100"; d2 <= "0011"; d3 <= "0011"; d4 <= "0000"; -- 334
    when "0000000101001111" => d1 <= "0101"; d2 <= "0011"; d3 <= "0011"; d4 <= "0000"; -- 335
    when "0000000101010000" => d1 <= "0110"; d2 <= "0011"; d3 <= "0011"; d4 <= "0000"; -- 336
    when "0000000101010001" => d1 <= "0111"; d2 <= "0011"; d3 <= "0011"; d4 <= "0000"; -- 337
    when "0000000101010010" => d1 <= "1000"; d2 <= "0011"; d3 <= "0011"; d4 <= "0000"; -- 338
    when "0000000101010011" => d1 <= "1001"; d2 <= "0011"; d3 <= "0011"; d4 <= "0000"; -- 339
    when "0000000101010100" => d1 <= "0000"; d2 <= "0100"; d3 <= "0011"; d4 <= "0000"; -- 340
    when "0000000101010101" => d1 <= "0001"; d2 <= "0100"; d3 <= "0011"; d4 <= "0000"; -- 341
    when "0000000101010110" => d1 <= "0010"; d2 <= "0100"; d3 <= "0011"; d4 <= "0000"; -- 342
    when "0000000101010111" => d1 <= "0011"; d2 <= "0100"; d3 <= "0011"; d4 <= "0000"; -- 343
    when "0000000101011000" => d1 <= "0100"; d2 <= "0100"; d3 <= "0011"; d4 <= "0000"; -- 344
    when "0000000101011001" => d1 <= "0101"; d2 <= "0100"; d3 <= "0011"; d4 <= "0000"; -- 345
    when "0000000101011010" => d1 <= "0110"; d2 <= "0100"; d3 <= "0011"; d4 <= "0000"; -- 346
    when "0000000101011011" => d1 <= "0111"; d2 <= "0100"; d3 <= "0011"; d4 <= "0000"; -- 347
    when "0000000101011100" => d1 <= "1000"; d2 <= "0100"; d3 <= "0011"; d4 <= "0000"; -- 348
    when "0000000101011101" => d1 <= "1001"; d2 <= "0100"; d3 <= "0011"; d4 <= "0000"; -- 349
    when "0000000101011110" => d1 <= "0000"; d2 <= "0101"; d3 <= "0011"; d4 <= "0000"; -- 350
    when "0000000101011111" => d1 <= "0001"; d2 <= "0101"; d3 <= "0011"; d4 <= "0000"; -- 351
    when "0000000101100000" => d1 <= "0010"; d2 <= "0101"; d3 <= "0011"; d4 <= "0000"; -- 352
    when "0000000101100001" => d1 <= "0011"; d2 <= "0101"; d3 <= "0011"; d4 <= "0000"; -- 353
    when "0000000101100010" => d1 <= "0100"; d2 <= "0101"; d3 <= "0011"; d4 <= "0000"; -- 354
    when "0000000101100011" => d1 <= "0101"; d2 <= "0101"; d3 <= "0011"; d4 <= "0000"; -- 355
    when "0000000101100100" => d1 <= "0110"; d2 <= "0101"; d3 <= "0011"; d4 <= "0000"; -- 356
    when "0000000101100101" => d1 <= "0111"; d2 <= "0101"; d3 <= "0011"; d4 <= "0000"; -- 357
    when "0000000101100110" => d1 <= "1000"; d2 <= "0101"; d3 <= "0011"; d4 <= "0000"; -- 358
    when "0000000101100111" => d1 <= "1001"; d2 <= "0101"; d3 <= "0011"; d4 <= "0000"; -- 359
    when "0000000101101000" => d1 <= "0000"; d2 <= "0110"; d3 <= "0011"; d4 <= "0000"; -- 360
    when "0000000101101001" => d1 <= "0001"; d2 <= "0110"; d3 <= "0011"; d4 <= "0000"; -- 361
    when "0000000101101010" => d1 <= "0010"; d2 <= "0110"; d3 <= "0011"; d4 <= "0000"; -- 362
    when "0000000101101011" => d1 <= "0011"; d2 <= "0110"; d3 <= "0011"; d4 <= "0000"; -- 363
    when "0000000101101100" => d1 <= "0100"; d2 <= "0110"; d3 <= "0011"; d4 <= "0000"; -- 364
    when "0000000101101101" => d1 <= "0101"; d2 <= "0110"; d3 <= "0011"; d4 <= "0000"; -- 365
    when "0000000101101110" => d1 <= "0110"; d2 <= "0110"; d3 <= "0011"; d4 <= "0000"; -- 366
    when "0000000101101111" => d1 <= "0111"; d2 <= "0110"; d3 <= "0011"; d4 <= "0000"; -- 367
    when "0000000101110000" => d1 <= "1000"; d2 <= "0110"; d3 <= "0011"; d4 <= "0000"; -- 368
    when "0000000101110001" => d1 <= "1001"; d2 <= "0110"; d3 <= "0011"; d4 <= "0000"; -- 369
    when "0000000101110010" => d1 <= "0000"; d2 <= "0111"; d3 <= "0011"; d4 <= "0000"; -- 370
    when "0000000101110011" => d1 <= "0001"; d2 <= "0111"; d3 <= "0011"; d4 <= "0000"; -- 371
    when "0000000101110100" => d1 <= "0010"; d2 <= "0111"; d3 <= "0011"; d4 <= "0000"; -- 372
    when "0000000101110101" => d1 <= "0011"; d2 <= "0111"; d3 <= "0011"; d4 <= "0000"; -- 373
    when "0000000101110110" => d1 <= "0100"; d2 <= "0111"; d3 <= "0011"; d4 <= "0000"; -- 374
    when "0000000101110111" => d1 <= "0101"; d2 <= "0111"; d3 <= "0011"; d4 <= "0000"; -- 375
    when "0000000101111000" => d1 <= "0110"; d2 <= "0111"; d3 <= "0011"; d4 <= "0000"; -- 376
    when "0000000101111001" => d1 <= "0111"; d2 <= "0111"; d3 <= "0011"; d4 <= "0000"; -- 377
    when "0000000101111010" => d1 <= "1000"; d2 <= "0111"; d3 <= "0011"; d4 <= "0000"; -- 378
    when "0000000101111011" => d1 <= "1001"; d2 <= "0111"; d3 <= "0011"; d4 <= "0000"; -- 379
    when "0000000101111100" => d1 <= "0000"; d2 <= "1000"; d3 <= "0011"; d4 <= "0000"; -- 380
    when "0000000101111101" => d1 <= "0001"; d2 <= "1000"; d3 <= "0011"; d4 <= "0000"; -- 381
    when "0000000101111110" => d1 <= "0010"; d2 <= "1000"; d3 <= "0011"; d4 <= "0000"; -- 382
    when "0000000101111111" => d1 <= "0011"; d2 <= "1000"; d3 <= "0011"; d4 <= "0000"; -- 383
    when "0000000110000000" => d1 <= "0100"; d2 <= "1000"; d3 <= "0011"; d4 <= "0000"; -- 384
    when "0000000110000001" => d1 <= "0101"; d2 <= "1000"; d3 <= "0011"; d4 <= "0000"; -- 385
    when "0000000110000010" => d1 <= "0110"; d2 <= "1000"; d3 <= "0011"; d4 <= "0000"; -- 386
    when "0000000110000011" => d1 <= "0111"; d2 <= "1000"; d3 <= "0011"; d4 <= "0000"; -- 387
    when "0000000110000100" => d1 <= "1000"; d2 <= "1000"; d3 <= "0011"; d4 <= "0000"; -- 388
    when "0000000110000101" => d1 <= "1001"; d2 <= "1000"; d3 <= "0011"; d4 <= "0000"; -- 389
    when "0000000110000110" => d1 <= "0000"; d2 <= "1001"; d3 <= "0011"; d4 <= "0000"; -- 390
    when "0000000110000111" => d1 <= "0001"; d2 <= "1001"; d3 <= "0011"; d4 <= "0000"; -- 391
    when "0000000110001000" => d1 <= "0010"; d2 <= "1001"; d3 <= "0011"; d4 <= "0000"; -- 392
    when "0000000110001001" => d1 <= "0011"; d2 <= "1001"; d3 <= "0011"; d4 <= "0000"; -- 393
    when "0000000110001010" => d1 <= "0100"; d2 <= "1001"; d3 <= "0011"; d4 <= "0000"; -- 394
    when "0000000110001011" => d1 <= "0101"; d2 <= "1001"; d3 <= "0011"; d4 <= "0000"; -- 395
    when "0000000110001100" => d1 <= "0110"; d2 <= "1001"; d3 <= "0011"; d4 <= "0000"; -- 396
    when "0000000110001101" => d1 <= "0111"; d2 <= "1001"; d3 <= "0011"; d4 <= "0000"; -- 397
    when "0000000110001110" => d1 <= "1000"; d2 <= "1001"; d3 <= "0011"; d4 <= "0000"; -- 398
    when "0000000110001111" => d1 <= "1001"; d2 <= "1001"; d3 <= "0011"; d4 <= "0000"; -- 399
    when "0000000110010000" => d1 <= "0000"; d2 <= "0000"; d3 <= "0100"; d4 <= "0000"; -- 400
    when "0000000110010001" => d1 <= "0001"; d2 <= "0000"; d3 <= "0100"; d4 <= "0000"; -- 401
    when "0000000110010010" => d1 <= "0010"; d2 <= "0000"; d3 <= "0100"; d4 <= "0000"; -- 402
    when "0000000110010011" => d1 <= "0011"; d2 <= "0000"; d3 <= "0100"; d4 <= "0000"; -- 403
    when "0000000110010100" => d1 <= "0100"; d2 <= "0000"; d3 <= "0100"; d4 <= "0000"; -- 404
    when "0000000110010101" => d1 <= "0101"; d2 <= "0000"; d3 <= "0100"; d4 <= "0000"; -- 405
    when "0000000110010110" => d1 <= "0110"; d2 <= "0000"; d3 <= "0100"; d4 <= "0000"; -- 406
    when "0000000110010111" => d1 <= "0111"; d2 <= "0000"; d3 <= "0100"; d4 <= "0000"; -- 407
    when "0000000110011000" => d1 <= "1000"; d2 <= "0000"; d3 <= "0100"; d4 <= "0000"; -- 408
    when "0000000110011001" => d1 <= "1001"; d2 <= "0000"; d3 <= "0100"; d4 <= "0000"; -- 409
    when "0000000110011010" => d1 <= "0000"; d2 <= "0001"; d3 <= "0100"; d4 <= "0000"; -- 410
    when "0000000110011011" => d1 <= "0001"; d2 <= "0001"; d3 <= "0100"; d4 <= "0000"; -- 411
    when "0000000110011100" => d1 <= "0010"; d2 <= "0001"; d3 <= "0100"; d4 <= "0000"; -- 412
    when "0000000110011101" => d1 <= "0011"; d2 <= "0001"; d3 <= "0100"; d4 <= "0000"; -- 413
    when "0000000110011110" => d1 <= "0100"; d2 <= "0001"; d3 <= "0100"; d4 <= "0000"; -- 414
    when "0000000110011111" => d1 <= "0101"; d2 <= "0001"; d3 <= "0100"; d4 <= "0000"; -- 415
    when "0000000110100000" => d1 <= "0110"; d2 <= "0001"; d3 <= "0100"; d4 <= "0000"; -- 416
    when "0000000110100001" => d1 <= "0111"; d2 <= "0001"; d3 <= "0100"; d4 <= "0000"; -- 417
    when "0000000110100010" => d1 <= "1000"; d2 <= "0001"; d3 <= "0100"; d4 <= "0000"; -- 418
    when "0000000110100011" => d1 <= "1001"; d2 <= "0001"; d3 <= "0100"; d4 <= "0000"; -- 419
    when "0000000110100100" => d1 <= "0000"; d2 <= "0010"; d3 <= "0100"; d4 <= "0000"; -- 420
    when "0000000110100101" => d1 <= "0001"; d2 <= "0010"; d3 <= "0100"; d4 <= "0000"; -- 421
    when "0000000110100110" => d1 <= "0010"; d2 <= "0010"; d3 <= "0100"; d4 <= "0000"; -- 422
    when "0000000110100111" => d1 <= "0011"; d2 <= "0010"; d3 <= "0100"; d4 <= "0000"; -- 423
    when "0000000110101000" => d1 <= "0100"; d2 <= "0010"; d3 <= "0100"; d4 <= "0000"; -- 424
    when "0000000110101001" => d1 <= "0101"; d2 <= "0010"; d3 <= "0100"; d4 <= "0000"; -- 425
    when "0000000110101010" => d1 <= "0110"; d2 <= "0010"; d3 <= "0100"; d4 <= "0000"; -- 426
    when "0000000110101011" => d1 <= "0111"; d2 <= "0010"; d3 <= "0100"; d4 <= "0000"; -- 427
    when "0000000110101100" => d1 <= "1000"; d2 <= "0010"; d3 <= "0100"; d4 <= "0000"; -- 428
    when "0000000110101101" => d1 <= "1001"; d2 <= "0010"; d3 <= "0100"; d4 <= "0000"; -- 429
    when "0000000110101110" => d1 <= "0000"; d2 <= "0011"; d3 <= "0100"; d4 <= "0000"; -- 430
    when "0000000110101111" => d1 <= "0001"; d2 <= "0011"; d3 <= "0100"; d4 <= "0000"; -- 431
    when "0000000110110000" => d1 <= "0010"; d2 <= "0011"; d3 <= "0100"; d4 <= "0000"; -- 432
    when "0000000110110001" => d1 <= "0011"; d2 <= "0011"; d3 <= "0100"; d4 <= "0000"; -- 433
    when "0000000110110010" => d1 <= "0100"; d2 <= "0011"; d3 <= "0100"; d4 <= "0000"; -- 434
    when "0000000110110011" => d1 <= "0101"; d2 <= "0011"; d3 <= "0100"; d4 <= "0000"; -- 435
    when "0000000110110100" => d1 <= "0110"; d2 <= "0011"; d3 <= "0100"; d4 <= "0000"; -- 436
    when "0000000110110101" => d1 <= "0111"; d2 <= "0011"; d3 <= "0100"; d4 <= "0000"; -- 437
    when "0000000110110110" => d1 <= "1000"; d2 <= "0011"; d3 <= "0100"; d4 <= "0000"; -- 438
    when "0000000110110111" => d1 <= "1001"; d2 <= "0011"; d3 <= "0100"; d4 <= "0000"; -- 439
    when "0000000110111000" => d1 <= "0000"; d2 <= "0100"; d3 <= "0100"; d4 <= "0000"; -- 440
    when "0000000110111001" => d1 <= "0001"; d2 <= "0100"; d3 <= "0100"; d4 <= "0000"; -- 441
    when "0000000110111010" => d1 <= "0010"; d2 <= "0100"; d3 <= "0100"; d4 <= "0000"; -- 442
    when "0000000110111011" => d1 <= "0011"; d2 <= "0100"; d3 <= "0100"; d4 <= "0000"; -- 443
    when "0000000110111100" => d1 <= "0100"; d2 <= "0100"; d3 <= "0100"; d4 <= "0000"; -- 444
    when "0000000110111101" => d1 <= "0101"; d2 <= "0100"; d3 <= "0100"; d4 <= "0000"; -- 445
    when "0000000110111110" => d1 <= "0110"; d2 <= "0100"; d3 <= "0100"; d4 <= "0000"; -- 446
    when "0000000110111111" => d1 <= "0111"; d2 <= "0100"; d3 <= "0100"; d4 <= "0000"; -- 447
    when "0000000111000000" => d1 <= "1000"; d2 <= "0100"; d3 <= "0100"; d4 <= "0000"; -- 448
    when "0000000111000001" => d1 <= "1001"; d2 <= "0100"; d3 <= "0100"; d4 <= "0000"; -- 449
    when "0000000111000010" => d1 <= "0000"; d2 <= "0101"; d3 <= "0100"; d4 <= "0000"; -- 450
    when "0000000111000011" => d1 <= "0001"; d2 <= "0101"; d3 <= "0100"; d4 <= "0000"; -- 451
    when "0000000111000100" => d1 <= "0010"; d2 <= "0101"; d3 <= "0100"; d4 <= "0000"; -- 452
    when "0000000111000101" => d1 <= "0011"; d2 <= "0101"; d3 <= "0100"; d4 <= "0000"; -- 453
    when "0000000111000110" => d1 <= "0100"; d2 <= "0101"; d3 <= "0100"; d4 <= "0000"; -- 454
    when "0000000111000111" => d1 <= "0101"; d2 <= "0101"; d3 <= "0100"; d4 <= "0000"; -- 455
    when "0000000111001000" => d1 <= "0110"; d2 <= "0101"; d3 <= "0100"; d4 <= "0000"; -- 456
    when "0000000111001001" => d1 <= "0111"; d2 <= "0101"; d3 <= "0100"; d4 <= "0000"; -- 457
    when "0000000111001010" => d1 <= "1000"; d2 <= "0101"; d3 <= "0100"; d4 <= "0000"; -- 458
    when "0000000111001011" => d1 <= "1001"; d2 <= "0101"; d3 <= "0100"; d4 <= "0000"; -- 459
    when "0000000111001100" => d1 <= "0000"; d2 <= "0110"; d3 <= "0100"; d4 <= "0000"; -- 460
    when "0000000111001101" => d1 <= "0001"; d2 <= "0110"; d3 <= "0100"; d4 <= "0000"; -- 461
    when "0000000111001110" => d1 <= "0010"; d2 <= "0110"; d3 <= "0100"; d4 <= "0000"; -- 462
    when "0000000111001111" => d1 <= "0011"; d2 <= "0110"; d3 <= "0100"; d4 <= "0000"; -- 463
    when "0000000111010000" => d1 <= "0100"; d2 <= "0110"; d3 <= "0100"; d4 <= "0000"; -- 464
    when "0000000111010001" => d1 <= "0101"; d2 <= "0110"; d3 <= "0100"; d4 <= "0000"; -- 465
    when "0000000111010010" => d1 <= "0110"; d2 <= "0110"; d3 <= "0100"; d4 <= "0000"; -- 466
    when "0000000111010011" => d1 <= "0111"; d2 <= "0110"; d3 <= "0100"; d4 <= "0000"; -- 467
    when "0000000111010100" => d1 <= "1000"; d2 <= "0110"; d3 <= "0100"; d4 <= "0000"; -- 468
    when "0000000111010101" => d1 <= "1001"; d2 <= "0110"; d3 <= "0100"; d4 <= "0000"; -- 469
    when "0000000111010110" => d1 <= "0000"; d2 <= "0111"; d3 <= "0100"; d4 <= "0000"; -- 470
    when "0000000111010111" => d1 <= "0001"; d2 <= "0111"; d3 <= "0100"; d4 <= "0000"; -- 471
    when "0000000111011000" => d1 <= "0010"; d2 <= "0111"; d3 <= "0100"; d4 <= "0000"; -- 472
    when "0000000111011001" => d1 <= "0011"; d2 <= "0111"; d3 <= "0100"; d4 <= "0000"; -- 473
    when "0000000111011010" => d1 <= "0100"; d2 <= "0111"; d3 <= "0100"; d4 <= "0000"; -- 474
    when "0000000111011011" => d1 <= "0101"; d2 <= "0111"; d3 <= "0100"; d4 <= "0000"; -- 475
    when "0000000111011100" => d1 <= "0110"; d2 <= "0111"; d3 <= "0100"; d4 <= "0000"; -- 476
    when "0000000111011101" => d1 <= "0111"; d2 <= "0111"; d3 <= "0100"; d4 <= "0000"; -- 477
    when "0000000111011110" => d1 <= "1000"; d2 <= "0111"; d3 <= "0100"; d4 <= "0000"; -- 478
    when "0000000111011111" => d1 <= "1001"; d2 <= "0111"; d3 <= "0100"; d4 <= "0000"; -- 479
    when "0000000111100000" => d1 <= "0000"; d2 <= "1000"; d3 <= "0100"; d4 <= "0000"; -- 480
    when "0000000111100001" => d1 <= "0001"; d2 <= "1000"; d3 <= "0100"; d4 <= "0000"; -- 481
    when "0000000111100010" => d1 <= "0010"; d2 <= "1000"; d3 <= "0100"; d4 <= "0000"; -- 482
    when "0000000111100011" => d1 <= "0011"; d2 <= "1000"; d3 <= "0100"; d4 <= "0000"; -- 483
    when "0000000111100100" => d1 <= "0100"; d2 <= "1000"; d3 <= "0100"; d4 <= "0000"; -- 484
    when "0000000111100101" => d1 <= "0101"; d2 <= "1000"; d3 <= "0100"; d4 <= "0000"; -- 485
    when "0000000111100110" => d1 <= "0110"; d2 <= "1000"; d3 <= "0100"; d4 <= "0000"; -- 486
    when "0000000111100111" => d1 <= "0111"; d2 <= "1000"; d3 <= "0100"; d4 <= "0000"; -- 487
    when "0000000111101000" => d1 <= "1000"; d2 <= "1000"; d3 <= "0100"; d4 <= "0000"; -- 488
    when "0000000111101001" => d1 <= "1001"; d2 <= "1000"; d3 <= "0100"; d4 <= "0000"; -- 489
    when "0000000111101010" => d1 <= "0000"; d2 <= "1001"; d3 <= "0100"; d4 <= "0000"; -- 490
    when "0000000111101011" => d1 <= "0001"; d2 <= "1001"; d3 <= "0100"; d4 <= "0000"; -- 491
    when "0000000111101100" => d1 <= "0010"; d2 <= "1001"; d3 <= "0100"; d4 <= "0000"; -- 492
    when "0000000111101101" => d1 <= "0011"; d2 <= "1001"; d3 <= "0100"; d4 <= "0000"; -- 493
    when "0000000111101110" => d1 <= "0100"; d2 <= "1001"; d3 <= "0100"; d4 <= "0000"; -- 494
    when "0000000111101111" => d1 <= "0101"; d2 <= "1001"; d3 <= "0100"; d4 <= "0000"; -- 495
    when "0000000111110000" => d1 <= "0110"; d2 <= "1001"; d3 <= "0100"; d4 <= "0000"; -- 496
    when "0000000111110001" => d1 <= "0111"; d2 <= "1001"; d3 <= "0100"; d4 <= "0000"; -- 497
    when "0000000111110010" => d1 <= "1000"; d2 <= "1001"; d3 <= "0100"; d4 <= "0000"; -- 498
    when "0000000111110011" => d1 <= "1001"; d2 <= "1001"; d3 <= "0100"; d4 <= "0000"; -- 499
    when "0000000111110100" => d1 <= "0000"; d2 <= "0000"; d3 <= "0101"; d4 <= "0000"; -- 500
    when "0000000111110101" => d1 <= "0001"; d2 <= "0000"; d3 <= "0101"; d4 <= "0000"; -- 501
    when "0000000111110110" => d1 <= "0010"; d2 <= "0000"; d3 <= "0101"; d4 <= "0000"; -- 502
    when "0000000111110111" => d1 <= "0011"; d2 <= "0000"; d3 <= "0101"; d4 <= "0000"; -- 503
    when "0000000111111000" => d1 <= "0100"; d2 <= "0000"; d3 <= "0101"; d4 <= "0000"; -- 504
    when "0000000111111001" => d1 <= "0101"; d2 <= "0000"; d3 <= "0101"; d4 <= "0000"; -- 505
    when "0000000111111010" => d1 <= "0110"; d2 <= "0000"; d3 <= "0101"; d4 <= "0000"; -- 506
    when "0000000111111011" => d1 <= "0111"; d2 <= "0000"; d3 <= "0101"; d4 <= "0000"; -- 507
    when "0000000111111100" => d1 <= "1000"; d2 <= "0000"; d3 <= "0101"; d4 <= "0000"; -- 508
    when "0000000111111101" => d1 <= "1001"; d2 <= "0000"; d3 <= "0101"; d4 <= "0000"; -- 509
    when "0000000111111110" => d1 <= "0000"; d2 <= "0001"; d3 <= "0101"; d4 <= "0000"; -- 510
    when "0000000111111111" => d1 <= "0001"; d2 <= "0001"; d3 <= "0101"; d4 <= "0000"; -- 511
    when "0000001000000000" => d1 <= "0010"; d2 <= "0001"; d3 <= "0101"; d4 <= "0000"; -- 512
    when "0000001000000001" => d1 <= "0011"; d2 <= "0001"; d3 <= "0101"; d4 <= "0000"; -- 513
    when "0000001000000010" => d1 <= "0100"; d2 <= "0001"; d3 <= "0101"; d4 <= "0000"; -- 514
    when "0000001000000011" => d1 <= "0101"; d2 <= "0001"; d3 <= "0101"; d4 <= "0000"; -- 515
    when "0000001000000100" => d1 <= "0110"; d2 <= "0001"; d3 <= "0101"; d4 <= "0000"; -- 516
    when "0000001000000101" => d1 <= "0111"; d2 <= "0001"; d3 <= "0101"; d4 <= "0000"; -- 517
    when "0000001000000110" => d1 <= "1000"; d2 <= "0001"; d3 <= "0101"; d4 <= "0000"; -- 518
    when "0000001000000111" => d1 <= "1001"; d2 <= "0001"; d3 <= "0101"; d4 <= "0000"; -- 519
    when "0000001000001000" => d1 <= "0000"; d2 <= "0010"; d3 <= "0101"; d4 <= "0000"; -- 520
    when "0000001000001001" => d1 <= "0001"; d2 <= "0010"; d3 <= "0101"; d4 <= "0000"; -- 521
    when "0000001000001010" => d1 <= "0010"; d2 <= "0010"; d3 <= "0101"; d4 <= "0000"; -- 522
    when "0000001000001011" => d1 <= "0011"; d2 <= "0010"; d3 <= "0101"; d4 <= "0000"; -- 523
    when "0000001000001100" => d1 <= "0100"; d2 <= "0010"; d3 <= "0101"; d4 <= "0000"; -- 524
    when "0000001000001101" => d1 <= "0101"; d2 <= "0010"; d3 <= "0101"; d4 <= "0000"; -- 525
    when "0000001000001110" => d1 <= "0110"; d2 <= "0010"; d3 <= "0101"; d4 <= "0000"; -- 526
    when "0000001000001111" => d1 <= "0111"; d2 <= "0010"; d3 <= "0101"; d4 <= "0000"; -- 527
    when "0000001000010000" => d1 <= "1000"; d2 <= "0010"; d3 <= "0101"; d4 <= "0000"; -- 528
    when "0000001000010001" => d1 <= "1001"; d2 <= "0010"; d3 <= "0101"; d4 <= "0000"; -- 529
    when "0000001000010010" => d1 <= "0000"; d2 <= "0011"; d3 <= "0101"; d4 <= "0000"; -- 530
    when "0000001000010011" => d1 <= "0001"; d2 <= "0011"; d3 <= "0101"; d4 <= "0000"; -- 531
    when "0000001000010100" => d1 <= "0010"; d2 <= "0011"; d3 <= "0101"; d4 <= "0000"; -- 532
    when "0000001000010101" => d1 <= "0011"; d2 <= "0011"; d3 <= "0101"; d4 <= "0000"; -- 533
    when "0000001000010110" => d1 <= "0100"; d2 <= "0011"; d3 <= "0101"; d4 <= "0000"; -- 534
    when "0000001000010111" => d1 <= "0101"; d2 <= "0011"; d3 <= "0101"; d4 <= "0000"; -- 535
    when "0000001000011000" => d1 <= "0110"; d2 <= "0011"; d3 <= "0101"; d4 <= "0000"; -- 536
    when "0000001000011001" => d1 <= "0111"; d2 <= "0011"; d3 <= "0101"; d4 <= "0000"; -- 537
    when "0000001000011010" => d1 <= "1000"; d2 <= "0011"; d3 <= "0101"; d4 <= "0000"; -- 538
    when "0000001000011011" => d1 <= "1001"; d2 <= "0011"; d3 <= "0101"; d4 <= "0000"; -- 539
    when "0000001000011100" => d1 <= "0000"; d2 <= "0100"; d3 <= "0101"; d4 <= "0000"; -- 540
    when "0000001000011101" => d1 <= "0001"; d2 <= "0100"; d3 <= "0101"; d4 <= "0000"; -- 541
    when "0000001000011110" => d1 <= "0010"; d2 <= "0100"; d3 <= "0101"; d4 <= "0000"; -- 542
    when "0000001000011111" => d1 <= "0011"; d2 <= "0100"; d3 <= "0101"; d4 <= "0000"; -- 543
    when "0000001000100000" => d1 <= "0100"; d2 <= "0100"; d3 <= "0101"; d4 <= "0000"; -- 544
    when "0000001000100001" => d1 <= "0101"; d2 <= "0100"; d3 <= "0101"; d4 <= "0000"; -- 545
    when "0000001000100010" => d1 <= "0110"; d2 <= "0100"; d3 <= "0101"; d4 <= "0000"; -- 546
    when "0000001000100011" => d1 <= "0111"; d2 <= "0100"; d3 <= "0101"; d4 <= "0000"; -- 547
    when "0000001000100100" => d1 <= "1000"; d2 <= "0100"; d3 <= "0101"; d4 <= "0000"; -- 548
    when "0000001000100101" => d1 <= "1001"; d2 <= "0100"; d3 <= "0101"; d4 <= "0000"; -- 549
    when "0000001000100110" => d1 <= "0000"; d2 <= "0101"; d3 <= "0101"; d4 <= "0000"; -- 550
    when "0000001000100111" => d1 <= "0001"; d2 <= "0101"; d3 <= "0101"; d4 <= "0000"; -- 551
    when "0000001000101000" => d1 <= "0010"; d2 <= "0101"; d3 <= "0101"; d4 <= "0000"; -- 552
    when "0000001000101001" => d1 <= "0011"; d2 <= "0101"; d3 <= "0101"; d4 <= "0000"; -- 553
    when "0000001000101010" => d1 <= "0100"; d2 <= "0101"; d3 <= "0101"; d4 <= "0000"; -- 554
    when "0000001000101011" => d1 <= "0101"; d2 <= "0101"; d3 <= "0101"; d4 <= "0000"; -- 555
    when "0000001000101100" => d1 <= "0110"; d2 <= "0101"; d3 <= "0101"; d4 <= "0000"; -- 556
    when "0000001000101101" => d1 <= "0111"; d2 <= "0101"; d3 <= "0101"; d4 <= "0000"; -- 557
    when "0000001000101110" => d1 <= "1000"; d2 <= "0101"; d3 <= "0101"; d4 <= "0000"; -- 558
    when "0000001000101111" => d1 <= "1001"; d2 <= "0101"; d3 <= "0101"; d4 <= "0000"; -- 559
    when "0000001000110000" => d1 <= "0000"; d2 <= "0110"; d3 <= "0101"; d4 <= "0000"; -- 560
    when "0000001000110001" => d1 <= "0001"; d2 <= "0110"; d3 <= "0101"; d4 <= "0000"; -- 561
    when "0000001000110010" => d1 <= "0010"; d2 <= "0110"; d3 <= "0101"; d4 <= "0000"; -- 562
    when "0000001000110011" => d1 <= "0011"; d2 <= "0110"; d3 <= "0101"; d4 <= "0000"; -- 563
    when "0000001000110100" => d1 <= "0100"; d2 <= "0110"; d3 <= "0101"; d4 <= "0000"; -- 564
    when "0000001000110101" => d1 <= "0101"; d2 <= "0110"; d3 <= "0101"; d4 <= "0000"; -- 565
    when "0000001000110110" => d1 <= "0110"; d2 <= "0110"; d3 <= "0101"; d4 <= "0000"; -- 566
    when "0000001000110111" => d1 <= "0111"; d2 <= "0110"; d3 <= "0101"; d4 <= "0000"; -- 567
    when "0000001000111000" => d1 <= "1000"; d2 <= "0110"; d3 <= "0101"; d4 <= "0000"; -- 568
    when "0000001000111001" => d1 <= "1001"; d2 <= "0110"; d3 <= "0101"; d4 <= "0000"; -- 569
    when "0000001000111010" => d1 <= "0000"; d2 <= "0111"; d3 <= "0101"; d4 <= "0000"; -- 570
    when "0000001000111011" => d1 <= "0001"; d2 <= "0111"; d3 <= "0101"; d4 <= "0000"; -- 571
    when "0000001000111100" => d1 <= "0010"; d2 <= "0111"; d3 <= "0101"; d4 <= "0000"; -- 572
    when "0000001000111101" => d1 <= "0011"; d2 <= "0111"; d3 <= "0101"; d4 <= "0000"; -- 573
    when "0000001000111110" => d1 <= "0100"; d2 <= "0111"; d3 <= "0101"; d4 <= "0000"; -- 574
    when "0000001000111111" => d1 <= "0101"; d2 <= "0111"; d3 <= "0101"; d4 <= "0000"; -- 575
    when "0000001001000000" => d1 <= "0110"; d2 <= "0111"; d3 <= "0101"; d4 <= "0000"; -- 576
    when "0000001001000001" => d1 <= "0111"; d2 <= "0111"; d3 <= "0101"; d4 <= "0000"; -- 577
    when "0000001001000010" => d1 <= "1000"; d2 <= "0111"; d3 <= "0101"; d4 <= "0000"; -- 578
    when "0000001001000011" => d1 <= "1001"; d2 <= "0111"; d3 <= "0101"; d4 <= "0000"; -- 579
    when "0000001001000100" => d1 <= "0000"; d2 <= "1000"; d3 <= "0101"; d4 <= "0000"; -- 580
    when "0000001001000101" => d1 <= "0001"; d2 <= "1000"; d3 <= "0101"; d4 <= "0000"; -- 581
    when "0000001001000110" => d1 <= "0010"; d2 <= "1000"; d3 <= "0101"; d4 <= "0000"; -- 582
    when "0000001001000111" => d1 <= "0011"; d2 <= "1000"; d3 <= "0101"; d4 <= "0000"; -- 583
    when "0000001001001000" => d1 <= "0100"; d2 <= "1000"; d3 <= "0101"; d4 <= "0000"; -- 584
    when "0000001001001001" => d1 <= "0101"; d2 <= "1000"; d3 <= "0101"; d4 <= "0000"; -- 585
    when "0000001001001010" => d1 <= "0110"; d2 <= "1000"; d3 <= "0101"; d4 <= "0000"; -- 586
    when "0000001001001011" => d1 <= "0111"; d2 <= "1000"; d3 <= "0101"; d4 <= "0000"; -- 587
    when "0000001001001100" => d1 <= "1000"; d2 <= "1000"; d3 <= "0101"; d4 <= "0000"; -- 588
    when "0000001001001101" => d1 <= "1001"; d2 <= "1000"; d3 <= "0101"; d4 <= "0000"; -- 589
    when "0000001001001110" => d1 <= "0000"; d2 <= "1001"; d3 <= "0101"; d4 <= "0000"; -- 590
    when "0000001001001111" => d1 <= "0001"; d2 <= "1001"; d3 <= "0101"; d4 <= "0000"; -- 591
    when "0000001001010000" => d1 <= "0010"; d2 <= "1001"; d3 <= "0101"; d4 <= "0000"; -- 592
    when "0000001001010001" => d1 <= "0011"; d2 <= "1001"; d3 <= "0101"; d4 <= "0000"; -- 593
    when "0000001001010010" => d1 <= "0100"; d2 <= "1001"; d3 <= "0101"; d4 <= "0000"; -- 594
    when "0000001001010011" => d1 <= "0101"; d2 <= "1001"; d3 <= "0101"; d4 <= "0000"; -- 595
    when "0000001001010100" => d1 <= "0110"; d2 <= "1001"; d3 <= "0101"; d4 <= "0000"; -- 596
    when "0000001001010101" => d1 <= "0111"; d2 <= "1001"; d3 <= "0101"; d4 <= "0000"; -- 597
    when "0000001001010110" => d1 <= "1000"; d2 <= "1001"; d3 <= "0101"; d4 <= "0000"; -- 598
    when "0000001001010111" => d1 <= "1001"; d2 <= "1001"; d3 <= "0101"; d4 <= "0000"; -- 599
    when "0000001001011000" => d1 <= "0000"; d2 <= "0000"; d3 <= "0110"; d4 <= "0000"; -- 600
    when "0000001001011001" => d1 <= "0001"; d2 <= "0000"; d3 <= "0110"; d4 <= "0000"; -- 601
    when "0000001001011010" => d1 <= "0010"; d2 <= "0000"; d3 <= "0110"; d4 <= "0000"; -- 602
    when "0000001001011011" => d1 <= "0011"; d2 <= "0000"; d3 <= "0110"; d4 <= "0000"; -- 603
    when "0000001001011100" => d1 <= "0100"; d2 <= "0000"; d3 <= "0110"; d4 <= "0000"; -- 604
    when "0000001001011101" => d1 <= "0101"; d2 <= "0000"; d3 <= "0110"; d4 <= "0000"; -- 605
    when "0000001001011110" => d1 <= "0110"; d2 <= "0000"; d3 <= "0110"; d4 <= "0000"; -- 606
    when "0000001001011111" => d1 <= "0111"; d2 <= "0000"; d3 <= "0110"; d4 <= "0000"; -- 607
    when "0000001001100000" => d1 <= "1000"; d2 <= "0000"; d3 <= "0110"; d4 <= "0000"; -- 608
    when "0000001001100001" => d1 <= "1001"; d2 <= "0000"; d3 <= "0110"; d4 <= "0000"; -- 609
    when "0000001001100010" => d1 <= "0000"; d2 <= "0001"; d3 <= "0110"; d4 <= "0000"; -- 610
    when "0000001001100011" => d1 <= "0001"; d2 <= "0001"; d3 <= "0110"; d4 <= "0000"; -- 611
    when "0000001001100100" => d1 <= "0010"; d2 <= "0001"; d3 <= "0110"; d4 <= "0000"; -- 612
    when "0000001001100101" => d1 <= "0011"; d2 <= "0001"; d3 <= "0110"; d4 <= "0000"; -- 613
    when "0000001001100110" => d1 <= "0100"; d2 <= "0001"; d3 <= "0110"; d4 <= "0000"; -- 614
    when "0000001001100111" => d1 <= "0101"; d2 <= "0001"; d3 <= "0110"; d4 <= "0000"; -- 615
    when "0000001001101000" => d1 <= "0110"; d2 <= "0001"; d3 <= "0110"; d4 <= "0000"; -- 616
    when "0000001001101001" => d1 <= "0111"; d2 <= "0001"; d3 <= "0110"; d4 <= "0000"; -- 617
    when "0000001001101010" => d1 <= "1000"; d2 <= "0001"; d3 <= "0110"; d4 <= "0000"; -- 618
    when "0000001001101011" => d1 <= "1001"; d2 <= "0001"; d3 <= "0110"; d4 <= "0000"; -- 619
    when "0000001001101100" => d1 <= "0000"; d2 <= "0010"; d3 <= "0110"; d4 <= "0000"; -- 620
    when "0000001001101101" => d1 <= "0001"; d2 <= "0010"; d3 <= "0110"; d4 <= "0000"; -- 621
    when "0000001001101110" => d1 <= "0010"; d2 <= "0010"; d3 <= "0110"; d4 <= "0000"; -- 622
    when "0000001001101111" => d1 <= "0011"; d2 <= "0010"; d3 <= "0110"; d4 <= "0000"; -- 623
    when "0000001001110000" => d1 <= "0100"; d2 <= "0010"; d3 <= "0110"; d4 <= "0000"; -- 624
    when "0000001001110001" => d1 <= "0101"; d2 <= "0010"; d3 <= "0110"; d4 <= "0000"; -- 625
    when "0000001001110010" => d1 <= "0110"; d2 <= "0010"; d3 <= "0110"; d4 <= "0000"; -- 626
    when "0000001001110011" => d1 <= "0111"; d2 <= "0010"; d3 <= "0110"; d4 <= "0000"; -- 627
    when "0000001001110100" => d1 <= "1000"; d2 <= "0010"; d3 <= "0110"; d4 <= "0000"; -- 628
    when "0000001001110101" => d1 <= "1001"; d2 <= "0010"; d3 <= "0110"; d4 <= "0000"; -- 629
    when "0000001001110110" => d1 <= "0000"; d2 <= "0011"; d3 <= "0110"; d4 <= "0000"; -- 630
    when "0000001001110111" => d1 <= "0001"; d2 <= "0011"; d3 <= "0110"; d4 <= "0000"; -- 631
    when "0000001001111000" => d1 <= "0010"; d2 <= "0011"; d3 <= "0110"; d4 <= "0000"; -- 632
    when "0000001001111001" => d1 <= "0011"; d2 <= "0011"; d3 <= "0110"; d4 <= "0000"; -- 633
    when "0000001001111010" => d1 <= "0100"; d2 <= "0011"; d3 <= "0110"; d4 <= "0000"; -- 634
    when "0000001001111011" => d1 <= "0101"; d2 <= "0011"; d3 <= "0110"; d4 <= "0000"; -- 635
    when "0000001001111100" => d1 <= "0110"; d2 <= "0011"; d3 <= "0110"; d4 <= "0000"; -- 636
    when "0000001001111101" => d1 <= "0111"; d2 <= "0011"; d3 <= "0110"; d4 <= "0000"; -- 637
    when "0000001001111110" => d1 <= "1000"; d2 <= "0011"; d3 <= "0110"; d4 <= "0000"; -- 638
    when "0000001001111111" => d1 <= "1001"; d2 <= "0011"; d3 <= "0110"; d4 <= "0000"; -- 639
    when "0000001010000000" => d1 <= "0000"; d2 <= "0100"; d3 <= "0110"; d4 <= "0000"; -- 640
    when "0000001010000001" => d1 <= "0001"; d2 <= "0100"; d3 <= "0110"; d4 <= "0000"; -- 641
    when "0000001010000010" => d1 <= "0010"; d2 <= "0100"; d3 <= "0110"; d4 <= "0000"; -- 642
    when "0000001010000011" => d1 <= "0011"; d2 <= "0100"; d3 <= "0110"; d4 <= "0000"; -- 643
    when "0000001010000100" => d1 <= "0100"; d2 <= "0100"; d3 <= "0110"; d4 <= "0000"; -- 644
    when "0000001010000101" => d1 <= "0101"; d2 <= "0100"; d3 <= "0110"; d4 <= "0000"; -- 645
    when "0000001010000110" => d1 <= "0110"; d2 <= "0100"; d3 <= "0110"; d4 <= "0000"; -- 646
    when "0000001010000111" => d1 <= "0111"; d2 <= "0100"; d3 <= "0110"; d4 <= "0000"; -- 647
    when "0000001010001000" => d1 <= "1000"; d2 <= "0100"; d3 <= "0110"; d4 <= "0000"; -- 648
    when "0000001010001001" => d1 <= "1001"; d2 <= "0100"; d3 <= "0110"; d4 <= "0000"; -- 649
    when "0000001010001010" => d1 <= "0000"; d2 <= "0101"; d3 <= "0110"; d4 <= "0000"; -- 650
    when "0000001010001011" => d1 <= "0001"; d2 <= "0101"; d3 <= "0110"; d4 <= "0000"; -- 651
    when "0000001010001100" => d1 <= "0010"; d2 <= "0101"; d3 <= "0110"; d4 <= "0000"; -- 652
    when "0000001010001101" => d1 <= "0011"; d2 <= "0101"; d3 <= "0110"; d4 <= "0000"; -- 653
    when "0000001010001110" => d1 <= "0100"; d2 <= "0101"; d3 <= "0110"; d4 <= "0000"; -- 654
    when "0000001010001111" => d1 <= "0101"; d2 <= "0101"; d3 <= "0110"; d4 <= "0000"; -- 655
    when "0000001010010000" => d1 <= "0110"; d2 <= "0101"; d3 <= "0110"; d4 <= "0000"; -- 656
    when "0000001010010001" => d1 <= "0111"; d2 <= "0101"; d3 <= "0110"; d4 <= "0000"; -- 657
    when "0000001010010010" => d1 <= "1000"; d2 <= "0101"; d3 <= "0110"; d4 <= "0000"; -- 658
    when "0000001010010011" => d1 <= "1001"; d2 <= "0101"; d3 <= "0110"; d4 <= "0000"; -- 659
    when "0000001010010100" => d1 <= "0000"; d2 <= "0110"; d3 <= "0110"; d4 <= "0000"; -- 660
    when "0000001010010101" => d1 <= "0001"; d2 <= "0110"; d3 <= "0110"; d4 <= "0000"; -- 661
    when "0000001010010110" => d1 <= "0010"; d2 <= "0110"; d3 <= "0110"; d4 <= "0000"; -- 662
    when "0000001010010111" => d1 <= "0011"; d2 <= "0110"; d3 <= "0110"; d4 <= "0000"; -- 663
    when "0000001010011000" => d1 <= "0100"; d2 <= "0110"; d3 <= "0110"; d4 <= "0000"; -- 664
    when "0000001010011001" => d1 <= "0101"; d2 <= "0110"; d3 <= "0110"; d4 <= "0000"; -- 665
    when "0000001010011010" => d1 <= "0110"; d2 <= "0110"; d3 <= "0110"; d4 <= "0000"; -- 666
    when "0000001010011011" => d1 <= "0111"; d2 <= "0110"; d3 <= "0110"; d4 <= "0000"; -- 667
    when "0000001010011100" => d1 <= "1000"; d2 <= "0110"; d3 <= "0110"; d4 <= "0000"; -- 668
    when "0000001010011101" => d1 <= "1001"; d2 <= "0110"; d3 <= "0110"; d4 <= "0000"; -- 669
    when "0000001010011110" => d1 <= "0000"; d2 <= "0111"; d3 <= "0110"; d4 <= "0000"; -- 670
    when "0000001010011111" => d1 <= "0001"; d2 <= "0111"; d3 <= "0110"; d4 <= "0000"; -- 671
    when "0000001010100000" => d1 <= "0010"; d2 <= "0111"; d3 <= "0110"; d4 <= "0000"; -- 672
    when "0000001010100001" => d1 <= "0011"; d2 <= "0111"; d3 <= "0110"; d4 <= "0000"; -- 673
    when "0000001010100010" => d1 <= "0100"; d2 <= "0111"; d3 <= "0110"; d4 <= "0000"; -- 674
    when "0000001010100011" => d1 <= "0101"; d2 <= "0111"; d3 <= "0110"; d4 <= "0000"; -- 675
    when "0000001010100100" => d1 <= "0110"; d2 <= "0111"; d3 <= "0110"; d4 <= "0000"; -- 676
    when "0000001010100101" => d1 <= "0111"; d2 <= "0111"; d3 <= "0110"; d4 <= "0000"; -- 677
    when "0000001010100110" => d1 <= "1000"; d2 <= "0111"; d3 <= "0110"; d4 <= "0000"; -- 678
    when "0000001010100111" => d1 <= "1001"; d2 <= "0111"; d3 <= "0110"; d4 <= "0000"; -- 679
    when "0000001010101000" => d1 <= "0000"; d2 <= "1000"; d3 <= "0110"; d4 <= "0000"; -- 680
    when "0000001010101001" => d1 <= "0001"; d2 <= "1000"; d3 <= "0110"; d4 <= "0000"; -- 681
    when "0000001010101010" => d1 <= "0010"; d2 <= "1000"; d3 <= "0110"; d4 <= "0000"; -- 682
    when "0000001010101011" => d1 <= "0011"; d2 <= "1000"; d3 <= "0110"; d4 <= "0000"; -- 683
    when "0000001010101100" => d1 <= "0100"; d2 <= "1000"; d3 <= "0110"; d4 <= "0000"; -- 684
    when "0000001010101101" => d1 <= "0101"; d2 <= "1000"; d3 <= "0110"; d4 <= "0000"; -- 685
    when "0000001010101110" => d1 <= "0110"; d2 <= "1000"; d3 <= "0110"; d4 <= "0000"; -- 686
    when "0000001010101111" => d1 <= "0111"; d2 <= "1000"; d3 <= "0110"; d4 <= "0000"; -- 687
    when "0000001010110000" => d1 <= "1000"; d2 <= "1000"; d3 <= "0110"; d4 <= "0000"; -- 688
    when "0000001010110001" => d1 <= "1001"; d2 <= "1000"; d3 <= "0110"; d4 <= "0000"; -- 689
    when "0000001010110010" => d1 <= "0000"; d2 <= "1001"; d3 <= "0110"; d4 <= "0000"; -- 690
    when "0000001010110011" => d1 <= "0001"; d2 <= "1001"; d3 <= "0110"; d4 <= "0000"; -- 691
    when "0000001010110100" => d1 <= "0010"; d2 <= "1001"; d3 <= "0110"; d4 <= "0000"; -- 692
    when "0000001010110101" => d1 <= "0011"; d2 <= "1001"; d3 <= "0110"; d4 <= "0000"; -- 693
    when "0000001010110110" => d1 <= "0100"; d2 <= "1001"; d3 <= "0110"; d4 <= "0000"; -- 694
    when "0000001010110111" => d1 <= "0101"; d2 <= "1001"; d3 <= "0110"; d4 <= "0000"; -- 695
    when "0000001010111000" => d1 <= "0110"; d2 <= "1001"; d3 <= "0110"; d4 <= "0000"; -- 696
    when "0000001010111001" => d1 <= "0111"; d2 <= "1001"; d3 <= "0110"; d4 <= "0000"; -- 697
    when "0000001010111010" => d1 <= "1000"; d2 <= "1001"; d3 <= "0110"; d4 <= "0000"; -- 698
    when "0000001010111011" => d1 <= "1001"; d2 <= "1001"; d3 <= "0110"; d4 <= "0000"; -- 699
    when "0000001010111100" => d1 <= "0000"; d2 <= "0000"; d3 <= "0111"; d4 <= "0000"; -- 700
    when "0000001010111101" => d1 <= "0001"; d2 <= "0000"; d3 <= "0111"; d4 <= "0000"; -- 701
    when "0000001010111110" => d1 <= "0010"; d2 <= "0000"; d3 <= "0111"; d4 <= "0000"; -- 702
    when "0000001010111111" => d1 <= "0011"; d2 <= "0000"; d3 <= "0111"; d4 <= "0000"; -- 703
    when "0000001011000000" => d1 <= "0100"; d2 <= "0000"; d3 <= "0111"; d4 <= "0000"; -- 704
    when "0000001011000001" => d1 <= "0101"; d2 <= "0000"; d3 <= "0111"; d4 <= "0000"; -- 705
    when "0000001011000010" => d1 <= "0110"; d2 <= "0000"; d3 <= "0111"; d4 <= "0000"; -- 706
    when "0000001011000011" => d1 <= "0111"; d2 <= "0000"; d3 <= "0111"; d4 <= "0000"; -- 707
    when "0000001011000100" => d1 <= "1000"; d2 <= "0000"; d3 <= "0111"; d4 <= "0000"; -- 708
    when "0000001011000101" => d1 <= "1001"; d2 <= "0000"; d3 <= "0111"; d4 <= "0000"; -- 709
    when "0000001011000110" => d1 <= "0000"; d2 <= "0001"; d3 <= "0111"; d4 <= "0000"; -- 710
    when "0000001011000111" => d1 <= "0001"; d2 <= "0001"; d3 <= "0111"; d4 <= "0000"; -- 711
    when "0000001011001000" => d1 <= "0010"; d2 <= "0001"; d3 <= "0111"; d4 <= "0000"; -- 712
    when "0000001011001001" => d1 <= "0011"; d2 <= "0001"; d3 <= "0111"; d4 <= "0000"; -- 713
    when "0000001011001010" => d1 <= "0100"; d2 <= "0001"; d3 <= "0111"; d4 <= "0000"; -- 714
    when "0000001011001011" => d1 <= "0101"; d2 <= "0001"; d3 <= "0111"; d4 <= "0000"; -- 715
    when "0000001011001100" => d1 <= "0110"; d2 <= "0001"; d3 <= "0111"; d4 <= "0000"; -- 716
    when "0000001011001101" => d1 <= "0111"; d2 <= "0001"; d3 <= "0111"; d4 <= "0000"; -- 717
    when "0000001011001110" => d1 <= "1000"; d2 <= "0001"; d3 <= "0111"; d4 <= "0000"; -- 718
    when "0000001011001111" => d1 <= "1001"; d2 <= "0001"; d3 <= "0111"; d4 <= "0000"; -- 719
    when "0000001011010000" => d1 <= "0000"; d2 <= "0010"; d3 <= "0111"; d4 <= "0000"; -- 720
    when "0000001011010001" => d1 <= "0001"; d2 <= "0010"; d3 <= "0111"; d4 <= "0000"; -- 721
    when "0000001011010010" => d1 <= "0010"; d2 <= "0010"; d3 <= "0111"; d4 <= "0000"; -- 722
    when "0000001011010011" => d1 <= "0011"; d2 <= "0010"; d3 <= "0111"; d4 <= "0000"; -- 723
    when "0000001011010100" => d1 <= "0100"; d2 <= "0010"; d3 <= "0111"; d4 <= "0000"; -- 724
    when "0000001011010101" => d1 <= "0101"; d2 <= "0010"; d3 <= "0111"; d4 <= "0000"; -- 725
    when "0000001011010110" => d1 <= "0110"; d2 <= "0010"; d3 <= "0111"; d4 <= "0000"; -- 726
    when "0000001011010111" => d1 <= "0111"; d2 <= "0010"; d3 <= "0111"; d4 <= "0000"; -- 727
    when "0000001011011000" => d1 <= "1000"; d2 <= "0010"; d3 <= "0111"; d4 <= "0000"; -- 728
    when "0000001011011001" => d1 <= "1001"; d2 <= "0010"; d3 <= "0111"; d4 <= "0000"; -- 729
    when "0000001011011010" => d1 <= "0000"; d2 <= "0011"; d3 <= "0111"; d4 <= "0000"; -- 730
    when "0000001011011011" => d1 <= "0001"; d2 <= "0011"; d3 <= "0111"; d4 <= "0000"; -- 731
    when "0000001011011100" => d1 <= "0010"; d2 <= "0011"; d3 <= "0111"; d4 <= "0000"; -- 732
    when "0000001011011101" => d1 <= "0011"; d2 <= "0011"; d3 <= "0111"; d4 <= "0000"; -- 733
    when "0000001011011110" => d1 <= "0100"; d2 <= "0011"; d3 <= "0111"; d4 <= "0000"; -- 734
    when "0000001011011111" => d1 <= "0101"; d2 <= "0011"; d3 <= "0111"; d4 <= "0000"; -- 735
    when "0000001011100000" => d1 <= "0110"; d2 <= "0011"; d3 <= "0111"; d4 <= "0000"; -- 736
    when "0000001011100001" => d1 <= "0111"; d2 <= "0011"; d3 <= "0111"; d4 <= "0000"; -- 737
    when "0000001011100010" => d1 <= "1000"; d2 <= "0011"; d3 <= "0111"; d4 <= "0000"; -- 738
    when "0000001011100011" => d1 <= "1001"; d2 <= "0011"; d3 <= "0111"; d4 <= "0000"; -- 739
    when "0000001011100100" => d1 <= "0000"; d2 <= "0100"; d3 <= "0111"; d4 <= "0000"; -- 740
    when "0000001011100101" => d1 <= "0001"; d2 <= "0100"; d3 <= "0111"; d4 <= "0000"; -- 741
    when "0000001011100110" => d1 <= "0010"; d2 <= "0100"; d3 <= "0111"; d4 <= "0000"; -- 742
    when "0000001011100111" => d1 <= "0011"; d2 <= "0100"; d3 <= "0111"; d4 <= "0000"; -- 743
    when "0000001011101000" => d1 <= "0100"; d2 <= "0100"; d3 <= "0111"; d4 <= "0000"; -- 744
    when "0000001011101001" => d1 <= "0101"; d2 <= "0100"; d3 <= "0111"; d4 <= "0000"; -- 745
    when "0000001011101010" => d1 <= "0110"; d2 <= "0100"; d3 <= "0111"; d4 <= "0000"; -- 746
    when "0000001011101011" => d1 <= "0111"; d2 <= "0100"; d3 <= "0111"; d4 <= "0000"; -- 747
    when "0000001011101100" => d1 <= "1000"; d2 <= "0100"; d3 <= "0111"; d4 <= "0000"; -- 748
    when "0000001011101101" => d1 <= "1001"; d2 <= "0100"; d3 <= "0111"; d4 <= "0000"; -- 749
    when "0000001011101110" => d1 <= "0000"; d2 <= "0101"; d3 <= "0111"; d4 <= "0000"; -- 750
    when "0000001011101111" => d1 <= "0001"; d2 <= "0101"; d3 <= "0111"; d4 <= "0000"; -- 751
    when "0000001011110000" => d1 <= "0010"; d2 <= "0101"; d3 <= "0111"; d4 <= "0000"; -- 752
    when "0000001011110001" => d1 <= "0011"; d2 <= "0101"; d3 <= "0111"; d4 <= "0000"; -- 753
    when "0000001011110010" => d1 <= "0100"; d2 <= "0101"; d3 <= "0111"; d4 <= "0000"; -- 754
    when "0000001011110011" => d1 <= "0101"; d2 <= "0101"; d3 <= "0111"; d4 <= "0000"; -- 755
    when "0000001011110100" => d1 <= "0110"; d2 <= "0101"; d3 <= "0111"; d4 <= "0000"; -- 756
    when "0000001011110101" => d1 <= "0111"; d2 <= "0101"; d3 <= "0111"; d4 <= "0000"; -- 757
    when "0000001011110110" => d1 <= "1000"; d2 <= "0101"; d3 <= "0111"; d4 <= "0000"; -- 758
    when "0000001011110111" => d1 <= "1001"; d2 <= "0101"; d3 <= "0111"; d4 <= "0000"; -- 759
    when "0000001011111000" => d1 <= "0000"; d2 <= "0110"; d3 <= "0111"; d4 <= "0000"; -- 760
    when "0000001011111001" => d1 <= "0001"; d2 <= "0110"; d3 <= "0111"; d4 <= "0000"; -- 761
    when "0000001011111010" => d1 <= "0010"; d2 <= "0110"; d3 <= "0111"; d4 <= "0000"; -- 762
    when "0000001011111011" => d1 <= "0011"; d2 <= "0110"; d3 <= "0111"; d4 <= "0000"; -- 763
    when "0000001011111100" => d1 <= "0100"; d2 <= "0110"; d3 <= "0111"; d4 <= "0000"; -- 764
    when "0000001011111101" => d1 <= "0101"; d2 <= "0110"; d3 <= "0111"; d4 <= "0000"; -- 765
    when "0000001011111110" => d1 <= "0110"; d2 <= "0110"; d3 <= "0111"; d4 <= "0000"; -- 766
    when "0000001011111111" => d1 <= "0111"; d2 <= "0110"; d3 <= "0111"; d4 <= "0000"; -- 767
    when "0000001100000000" => d1 <= "1000"; d2 <= "0110"; d3 <= "0111"; d4 <= "0000"; -- 768
    when "0000001100000001" => d1 <= "1001"; d2 <= "0110"; d3 <= "0111"; d4 <= "0000"; -- 769
    when "0000001100000010" => d1 <= "0000"; d2 <= "0111"; d3 <= "0111"; d4 <= "0000"; -- 770
    when "0000001100000011" => d1 <= "0001"; d2 <= "0111"; d3 <= "0111"; d4 <= "0000"; -- 771
    when "0000001100000100" => d1 <= "0010"; d2 <= "0111"; d3 <= "0111"; d4 <= "0000"; -- 772
    when "0000001100000101" => d1 <= "0011"; d2 <= "0111"; d3 <= "0111"; d4 <= "0000"; -- 773
    when "0000001100000110" => d1 <= "0100"; d2 <= "0111"; d3 <= "0111"; d4 <= "0000"; -- 774
    when "0000001100000111" => d1 <= "0101"; d2 <= "0111"; d3 <= "0111"; d4 <= "0000"; -- 775
    when "0000001100001000" => d1 <= "0110"; d2 <= "0111"; d3 <= "0111"; d4 <= "0000"; -- 776
    when "0000001100001001" => d1 <= "0111"; d2 <= "0111"; d3 <= "0111"; d4 <= "0000"; -- 777
    when "0000001100001010" => d1 <= "1000"; d2 <= "0111"; d3 <= "0111"; d4 <= "0000"; -- 778
    when "0000001100001011" => d1 <= "1001"; d2 <= "0111"; d3 <= "0111"; d4 <= "0000"; -- 779
    when "0000001100001100" => d1 <= "0000"; d2 <= "1000"; d3 <= "0111"; d4 <= "0000"; -- 780
    when "0000001100001101" => d1 <= "0001"; d2 <= "1000"; d3 <= "0111"; d4 <= "0000"; -- 781
    when "0000001100001110" => d1 <= "0010"; d2 <= "1000"; d3 <= "0111"; d4 <= "0000"; -- 782
    when "0000001100001111" => d1 <= "0011"; d2 <= "1000"; d3 <= "0111"; d4 <= "0000"; -- 783
    when "0000001100010000" => d1 <= "0100"; d2 <= "1000"; d3 <= "0111"; d4 <= "0000"; -- 784
    when "0000001100010001" => d1 <= "0101"; d2 <= "1000"; d3 <= "0111"; d4 <= "0000"; -- 785
    when "0000001100010010" => d1 <= "0110"; d2 <= "1000"; d3 <= "0111"; d4 <= "0000"; -- 786
    when "0000001100010011" => d1 <= "0111"; d2 <= "1000"; d3 <= "0111"; d4 <= "0000"; -- 787
    when "0000001100010100" => d1 <= "1000"; d2 <= "1000"; d3 <= "0111"; d4 <= "0000"; -- 788
    when "0000001100010101" => d1 <= "1001"; d2 <= "1000"; d3 <= "0111"; d4 <= "0000"; -- 789
    when "0000001100010110" => d1 <= "0000"; d2 <= "1001"; d3 <= "0111"; d4 <= "0000"; -- 790
    when "0000001100010111" => d1 <= "0001"; d2 <= "1001"; d3 <= "0111"; d4 <= "0000"; -- 791
    when "0000001100011000" => d1 <= "0010"; d2 <= "1001"; d3 <= "0111"; d4 <= "0000"; -- 792
    when "0000001100011001" => d1 <= "0011"; d2 <= "1001"; d3 <= "0111"; d4 <= "0000"; -- 793
    when "0000001100011010" => d1 <= "0100"; d2 <= "1001"; d3 <= "0111"; d4 <= "0000"; -- 794
    when "0000001100011011" => d1 <= "0101"; d2 <= "1001"; d3 <= "0111"; d4 <= "0000"; -- 795
    when "0000001100011100" => d1 <= "0110"; d2 <= "1001"; d3 <= "0111"; d4 <= "0000"; -- 796
    when "0000001100011101" => d1 <= "0111"; d2 <= "1001"; d3 <= "0111"; d4 <= "0000"; -- 797
    when "0000001100011110" => d1 <= "1000"; d2 <= "1001"; d3 <= "0111"; d4 <= "0000"; -- 798
    when "0000001100011111" => d1 <= "1001"; d2 <= "1001"; d3 <= "0111"; d4 <= "0000"; -- 799
    when "0000001100100000" => d1 <= "0000"; d2 <= "0000"; d3 <= "1000"; d4 <= "0000"; -- 800
    when "0000001100100001" => d1 <= "0001"; d2 <= "0000"; d3 <= "1000"; d4 <= "0000"; -- 801
    when "0000001100100010" => d1 <= "0010"; d2 <= "0000"; d3 <= "1000"; d4 <= "0000"; -- 802
    when "0000001100100011" => d1 <= "0011"; d2 <= "0000"; d3 <= "1000"; d4 <= "0000"; -- 803
    when "0000001100100100" => d1 <= "0100"; d2 <= "0000"; d3 <= "1000"; d4 <= "0000"; -- 804
    when "0000001100100101" => d1 <= "0101"; d2 <= "0000"; d3 <= "1000"; d4 <= "0000"; -- 805
    when "0000001100100110" => d1 <= "0110"; d2 <= "0000"; d3 <= "1000"; d4 <= "0000"; -- 806
    when "0000001100100111" => d1 <= "0111"; d2 <= "0000"; d3 <= "1000"; d4 <= "0000"; -- 807
    when "0000001100101000" => d1 <= "1000"; d2 <= "0000"; d3 <= "1000"; d4 <= "0000"; -- 808
    when "0000001100101001" => d1 <= "1001"; d2 <= "0000"; d3 <= "1000"; d4 <= "0000"; -- 809
    when "0000001100101010" => d1 <= "0000"; d2 <= "0001"; d3 <= "1000"; d4 <= "0000"; -- 810
    when "0000001100101011" => d1 <= "0001"; d2 <= "0001"; d3 <= "1000"; d4 <= "0000"; -- 811
    when "0000001100101100" => d1 <= "0010"; d2 <= "0001"; d3 <= "1000"; d4 <= "0000"; -- 812
    when "0000001100101101" => d1 <= "0011"; d2 <= "0001"; d3 <= "1000"; d4 <= "0000"; -- 813
    when "0000001100101110" => d1 <= "0100"; d2 <= "0001"; d3 <= "1000"; d4 <= "0000"; -- 814
    when "0000001100101111" => d1 <= "0101"; d2 <= "0001"; d3 <= "1000"; d4 <= "0000"; -- 815
    when "0000001100110000" => d1 <= "0110"; d2 <= "0001"; d3 <= "1000"; d4 <= "0000"; -- 816
    when "0000001100110001" => d1 <= "0111"; d2 <= "0001"; d3 <= "1000"; d4 <= "0000"; -- 817
    when "0000001100110010" => d1 <= "1000"; d2 <= "0001"; d3 <= "1000"; d4 <= "0000"; -- 818
    when "0000001100110011" => d1 <= "1001"; d2 <= "0001"; d3 <= "1000"; d4 <= "0000"; -- 819
    when "0000001100110100" => d1 <= "0000"; d2 <= "0010"; d3 <= "1000"; d4 <= "0000"; -- 820
    when "0000001100110101" => d1 <= "0001"; d2 <= "0010"; d3 <= "1000"; d4 <= "0000"; -- 821
    when "0000001100110110" => d1 <= "0010"; d2 <= "0010"; d3 <= "1000"; d4 <= "0000"; -- 822
    when "0000001100110111" => d1 <= "0011"; d2 <= "0010"; d3 <= "1000"; d4 <= "0000"; -- 823
    when "0000001100111000" => d1 <= "0100"; d2 <= "0010"; d3 <= "1000"; d4 <= "0000"; -- 824
    when "0000001100111001" => d1 <= "0101"; d2 <= "0010"; d3 <= "1000"; d4 <= "0000"; -- 825
    when "0000001100111010" => d1 <= "0110"; d2 <= "0010"; d3 <= "1000"; d4 <= "0000"; -- 826
    when "0000001100111011" => d1 <= "0111"; d2 <= "0010"; d3 <= "1000"; d4 <= "0000"; -- 827
    when "0000001100111100" => d1 <= "1000"; d2 <= "0010"; d3 <= "1000"; d4 <= "0000"; -- 828
    when "0000001100111101" => d1 <= "1001"; d2 <= "0010"; d3 <= "1000"; d4 <= "0000"; -- 829
    when "0000001100111110" => d1 <= "0000"; d2 <= "0011"; d3 <= "1000"; d4 <= "0000"; -- 830
    when "0000001100111111" => d1 <= "0001"; d2 <= "0011"; d3 <= "1000"; d4 <= "0000"; -- 831
    when "0000001101000000" => d1 <= "0010"; d2 <= "0011"; d3 <= "1000"; d4 <= "0000"; -- 832
    when "0000001101000001" => d1 <= "0011"; d2 <= "0011"; d3 <= "1000"; d4 <= "0000"; -- 833
    when "0000001101000010" => d1 <= "0100"; d2 <= "0011"; d3 <= "1000"; d4 <= "0000"; -- 834
    when "0000001101000011" => d1 <= "0101"; d2 <= "0011"; d3 <= "1000"; d4 <= "0000"; -- 835
    when "0000001101000100" => d1 <= "0110"; d2 <= "0011"; d3 <= "1000"; d4 <= "0000"; -- 836
    when "0000001101000101" => d1 <= "0111"; d2 <= "0011"; d3 <= "1000"; d4 <= "0000"; -- 837
    when "0000001101000110" => d1 <= "1000"; d2 <= "0011"; d3 <= "1000"; d4 <= "0000"; -- 838
    when "0000001101000111" => d1 <= "1001"; d2 <= "0011"; d3 <= "1000"; d4 <= "0000"; -- 839
    when "0000001101001000" => d1 <= "0000"; d2 <= "0100"; d3 <= "1000"; d4 <= "0000"; -- 840
    when "0000001101001001" => d1 <= "0001"; d2 <= "0100"; d3 <= "1000"; d4 <= "0000"; -- 841
    when "0000001101001010" => d1 <= "0010"; d2 <= "0100"; d3 <= "1000"; d4 <= "0000"; -- 842
    when "0000001101001011" => d1 <= "0011"; d2 <= "0100"; d3 <= "1000"; d4 <= "0000"; -- 843
    when "0000001101001100" => d1 <= "0100"; d2 <= "0100"; d3 <= "1000"; d4 <= "0000"; -- 844
    when "0000001101001101" => d1 <= "0101"; d2 <= "0100"; d3 <= "1000"; d4 <= "0000"; -- 845
    when "0000001101001110" => d1 <= "0110"; d2 <= "0100"; d3 <= "1000"; d4 <= "0000"; -- 846
    when "0000001101001111" => d1 <= "0111"; d2 <= "0100"; d3 <= "1000"; d4 <= "0000"; -- 847
    when "0000001101010000" => d1 <= "1000"; d2 <= "0100"; d3 <= "1000"; d4 <= "0000"; -- 848
    when "0000001101010001" => d1 <= "1001"; d2 <= "0100"; d3 <= "1000"; d4 <= "0000"; -- 849
    when "0000001101010010" => d1 <= "0000"; d2 <= "0101"; d3 <= "1000"; d4 <= "0000"; -- 850
    when "0000001101010011" => d1 <= "0001"; d2 <= "0101"; d3 <= "1000"; d4 <= "0000"; -- 851
    when "0000001101010100" => d1 <= "0010"; d2 <= "0101"; d3 <= "1000"; d4 <= "0000"; -- 852
    when "0000001101010101" => d1 <= "0011"; d2 <= "0101"; d3 <= "1000"; d4 <= "0000"; -- 853
    when "0000001101010110" => d1 <= "0100"; d2 <= "0101"; d3 <= "1000"; d4 <= "0000"; -- 854
    when "0000001101010111" => d1 <= "0101"; d2 <= "0101"; d3 <= "1000"; d4 <= "0000"; -- 855
    when "0000001101011000" => d1 <= "0110"; d2 <= "0101"; d3 <= "1000"; d4 <= "0000"; -- 856
    when "0000001101011001" => d1 <= "0111"; d2 <= "0101"; d3 <= "1000"; d4 <= "0000"; -- 857
    when "0000001101011010" => d1 <= "1000"; d2 <= "0101"; d3 <= "1000"; d4 <= "0000"; -- 858
    when "0000001101011011" => d1 <= "1001"; d2 <= "0101"; d3 <= "1000"; d4 <= "0000"; -- 859
    when "0000001101011100" => d1 <= "0000"; d2 <= "0110"; d3 <= "1000"; d4 <= "0000"; -- 860
    when "0000001101011101" => d1 <= "0001"; d2 <= "0110"; d3 <= "1000"; d4 <= "0000"; -- 861
    when "0000001101011110" => d1 <= "0010"; d2 <= "0110"; d3 <= "1000"; d4 <= "0000"; -- 862
    when "0000001101011111" => d1 <= "0011"; d2 <= "0110"; d3 <= "1000"; d4 <= "0000"; -- 863
    when "0000001101100000" => d1 <= "0100"; d2 <= "0110"; d3 <= "1000"; d4 <= "0000"; -- 864
    when "0000001101100001" => d1 <= "0101"; d2 <= "0110"; d3 <= "1000"; d4 <= "0000"; -- 865
    when "0000001101100010" => d1 <= "0110"; d2 <= "0110"; d3 <= "1000"; d4 <= "0000"; -- 866
    when "0000001101100011" => d1 <= "0111"; d2 <= "0110"; d3 <= "1000"; d4 <= "0000"; -- 867
    when "0000001101100100" => d1 <= "1000"; d2 <= "0110"; d3 <= "1000"; d4 <= "0000"; -- 868
    when "0000001101100101" => d1 <= "1001"; d2 <= "0110"; d3 <= "1000"; d4 <= "0000"; -- 869
    when "0000001101100110" => d1 <= "0000"; d2 <= "0111"; d3 <= "1000"; d4 <= "0000"; -- 870
    when "0000001101100111" => d1 <= "0001"; d2 <= "0111"; d3 <= "1000"; d4 <= "0000"; -- 871
    when "0000001101101000" => d1 <= "0010"; d2 <= "0111"; d3 <= "1000"; d4 <= "0000"; -- 872
    when "0000001101101001" => d1 <= "0011"; d2 <= "0111"; d3 <= "1000"; d4 <= "0000"; -- 873
    when "0000001101101010" => d1 <= "0100"; d2 <= "0111"; d3 <= "1000"; d4 <= "0000"; -- 874
    when "0000001101101011" => d1 <= "0101"; d2 <= "0111"; d3 <= "1000"; d4 <= "0000"; -- 875
    when "0000001101101100" => d1 <= "0110"; d2 <= "0111"; d3 <= "1000"; d4 <= "0000"; -- 876
    when "0000001101101101" => d1 <= "0111"; d2 <= "0111"; d3 <= "1000"; d4 <= "0000"; -- 877
    when "0000001101101110" => d1 <= "1000"; d2 <= "0111"; d3 <= "1000"; d4 <= "0000"; -- 878
    when "0000001101101111" => d1 <= "1001"; d2 <= "0111"; d3 <= "1000"; d4 <= "0000"; -- 879
    when "0000001101110000" => d1 <= "0000"; d2 <= "1000"; d3 <= "1000"; d4 <= "0000"; -- 880
    when "0000001101110001" => d1 <= "0001"; d2 <= "1000"; d3 <= "1000"; d4 <= "0000"; -- 881
    when "0000001101110010" => d1 <= "0010"; d2 <= "1000"; d3 <= "1000"; d4 <= "0000"; -- 882
    when "0000001101110011" => d1 <= "0011"; d2 <= "1000"; d3 <= "1000"; d4 <= "0000"; -- 883
    when "0000001101110100" => d1 <= "0100"; d2 <= "1000"; d3 <= "1000"; d4 <= "0000"; -- 884
    when "0000001101110101" => d1 <= "0101"; d2 <= "1000"; d3 <= "1000"; d4 <= "0000"; -- 885
    when "0000001101110110" => d1 <= "0110"; d2 <= "1000"; d3 <= "1000"; d4 <= "0000"; -- 886
    when "0000001101110111" => d1 <= "0111"; d2 <= "1000"; d3 <= "1000"; d4 <= "0000"; -- 887
    when "0000001101111000" => d1 <= "1000"; d2 <= "1000"; d3 <= "1000"; d4 <= "0000"; -- 888
    when "0000001101111001" => d1 <= "1001"; d2 <= "1000"; d3 <= "1000"; d4 <= "0000"; -- 889
    when "0000001101111010" => d1 <= "0000"; d2 <= "1001"; d3 <= "1000"; d4 <= "0000"; -- 890
    when "0000001101111011" => d1 <= "0001"; d2 <= "1001"; d3 <= "1000"; d4 <= "0000"; -- 891
    when "0000001101111100" => d1 <= "0010"; d2 <= "1001"; d3 <= "1000"; d4 <= "0000"; -- 892
    when "0000001101111101" => d1 <= "0011"; d2 <= "1001"; d3 <= "1000"; d4 <= "0000"; -- 893
    when "0000001101111110" => d1 <= "0100"; d2 <= "1001"; d3 <= "1000"; d4 <= "0000"; -- 894
    when "0000001101111111" => d1 <= "0101"; d2 <= "1001"; d3 <= "1000"; d4 <= "0000"; -- 895
    when "0000001110000000" => d1 <= "0110"; d2 <= "1001"; d3 <= "1000"; d4 <= "0000"; -- 896
    when "0000001110000001" => d1 <= "0111"; d2 <= "1001"; d3 <= "1000"; d4 <= "0000"; -- 897
    when "0000001110000010" => d1 <= "1000"; d2 <= "1001"; d3 <= "1000"; d4 <= "0000"; -- 898
    when "0000001110000011" => d1 <= "1001"; d2 <= "1001"; d3 <= "1000"; d4 <= "0000"; -- 899
    when "0000001110000100" => d1 <= "0000"; d2 <= "0000"; d3 <= "1001"; d4 <= "0000"; -- 900
    when "0000001110000101" => d1 <= "0001"; d2 <= "0000"; d3 <= "1001"; d4 <= "0000"; -- 901
    when "0000001110000110" => d1 <= "0010"; d2 <= "0000"; d3 <= "1001"; d4 <= "0000"; -- 902
    when "0000001110000111" => d1 <= "0011"; d2 <= "0000"; d3 <= "1001"; d4 <= "0000"; -- 903
    when "0000001110001000" => d1 <= "0100"; d2 <= "0000"; d3 <= "1001"; d4 <= "0000"; -- 904
    when "0000001110001001" => d1 <= "0101"; d2 <= "0000"; d3 <= "1001"; d4 <= "0000"; -- 905
    when "0000001110001010" => d1 <= "0110"; d2 <= "0000"; d3 <= "1001"; d4 <= "0000"; -- 906
    when "0000001110001011" => d1 <= "0111"; d2 <= "0000"; d3 <= "1001"; d4 <= "0000"; -- 907
    when "0000001110001100" => d1 <= "1000"; d2 <= "0000"; d3 <= "1001"; d4 <= "0000"; -- 908
    when "0000001110001101" => d1 <= "1001"; d2 <= "0000"; d3 <= "1001"; d4 <= "0000"; -- 909
    when "0000001110001110" => d1 <= "0000"; d2 <= "0001"; d3 <= "1001"; d4 <= "0000"; -- 910
    when "0000001110001111" => d1 <= "0001"; d2 <= "0001"; d3 <= "1001"; d4 <= "0000"; -- 911
    when "0000001110010000" => d1 <= "0010"; d2 <= "0001"; d3 <= "1001"; d4 <= "0000"; -- 912
    when "0000001110010001" => d1 <= "0011"; d2 <= "0001"; d3 <= "1001"; d4 <= "0000"; -- 913
    when "0000001110010010" => d1 <= "0100"; d2 <= "0001"; d3 <= "1001"; d4 <= "0000"; -- 914
    when "0000001110010011" => d1 <= "0101"; d2 <= "0001"; d3 <= "1001"; d4 <= "0000"; -- 915
    when "0000001110010100" => d1 <= "0110"; d2 <= "0001"; d3 <= "1001"; d4 <= "0000"; -- 916
    when "0000001110010101" => d1 <= "0111"; d2 <= "0001"; d3 <= "1001"; d4 <= "0000"; -- 917
    when "0000001110010110" => d1 <= "1000"; d2 <= "0001"; d3 <= "1001"; d4 <= "0000"; -- 918
    when "0000001110010111" => d1 <= "1001"; d2 <= "0001"; d3 <= "1001"; d4 <= "0000"; -- 919
    when "0000001110011000" => d1 <= "0000"; d2 <= "0010"; d3 <= "1001"; d4 <= "0000"; -- 920
    when "0000001110011001" => d1 <= "0001"; d2 <= "0010"; d3 <= "1001"; d4 <= "0000"; -- 921
    when "0000001110011010" => d1 <= "0010"; d2 <= "0010"; d3 <= "1001"; d4 <= "0000"; -- 922
    when "0000001110011011" => d1 <= "0011"; d2 <= "0010"; d3 <= "1001"; d4 <= "0000"; -- 923
    when "0000001110011100" => d1 <= "0100"; d2 <= "0010"; d3 <= "1001"; d4 <= "0000"; -- 924
    when "0000001110011101" => d1 <= "0101"; d2 <= "0010"; d3 <= "1001"; d4 <= "0000"; -- 925
    when "0000001110011110" => d1 <= "0110"; d2 <= "0010"; d3 <= "1001"; d4 <= "0000"; -- 926
    when "0000001110011111" => d1 <= "0111"; d2 <= "0010"; d3 <= "1001"; d4 <= "0000"; -- 927
    when "0000001110100000" => d1 <= "1000"; d2 <= "0010"; d3 <= "1001"; d4 <= "0000"; -- 928
    when "0000001110100001" => d1 <= "1001"; d2 <= "0010"; d3 <= "1001"; d4 <= "0000"; -- 929
    when "0000001110100010" => d1 <= "0000"; d2 <= "0011"; d3 <= "1001"; d4 <= "0000"; -- 930
    when "0000001110100011" => d1 <= "0001"; d2 <= "0011"; d3 <= "1001"; d4 <= "0000"; -- 931
    when "0000001110100100" => d1 <= "0010"; d2 <= "0011"; d3 <= "1001"; d4 <= "0000"; -- 932
    when "0000001110100101" => d1 <= "0011"; d2 <= "0011"; d3 <= "1001"; d4 <= "0000"; -- 933
    when "0000001110100110" => d1 <= "0100"; d2 <= "0011"; d3 <= "1001"; d4 <= "0000"; -- 934
    when "0000001110100111" => d1 <= "0101"; d2 <= "0011"; d3 <= "1001"; d4 <= "0000"; -- 935
    when "0000001110101000" => d1 <= "0110"; d2 <= "0011"; d3 <= "1001"; d4 <= "0000"; -- 936
    when "0000001110101001" => d1 <= "0111"; d2 <= "0011"; d3 <= "1001"; d4 <= "0000"; -- 937
    when "0000001110101010" => d1 <= "1000"; d2 <= "0011"; d3 <= "1001"; d4 <= "0000"; -- 938
    when "0000001110101011" => d1 <= "1001"; d2 <= "0011"; d3 <= "1001"; d4 <= "0000"; -- 939
    when "0000001110101100" => d1 <= "0000"; d2 <= "0100"; d3 <= "1001"; d4 <= "0000"; -- 940
    when "0000001110101101" => d1 <= "0001"; d2 <= "0100"; d3 <= "1001"; d4 <= "0000"; -- 941
    when "0000001110101110" => d1 <= "0010"; d2 <= "0100"; d3 <= "1001"; d4 <= "0000"; -- 942
    when "0000001110101111" => d1 <= "0011"; d2 <= "0100"; d3 <= "1001"; d4 <= "0000"; -- 943
    when "0000001110110000" => d1 <= "0100"; d2 <= "0100"; d3 <= "1001"; d4 <= "0000"; -- 944
    when "0000001110110001" => d1 <= "0101"; d2 <= "0100"; d3 <= "1001"; d4 <= "0000"; -- 945
    when "0000001110110010" => d1 <= "0110"; d2 <= "0100"; d3 <= "1001"; d4 <= "0000"; -- 946
    when "0000001110110011" => d1 <= "0111"; d2 <= "0100"; d3 <= "1001"; d4 <= "0000"; -- 947
    when "0000001110110100" => d1 <= "1000"; d2 <= "0100"; d3 <= "1001"; d4 <= "0000"; -- 948
    when "0000001110110101" => d1 <= "1001"; d2 <= "0100"; d3 <= "1001"; d4 <= "0000"; -- 949
    when "0000001110110110" => d1 <= "0000"; d2 <= "0101"; d3 <= "1001"; d4 <= "0000"; -- 950
    when "0000001110110111" => d1 <= "0001"; d2 <= "0101"; d3 <= "1001"; d4 <= "0000"; -- 951
    when "0000001110111000" => d1 <= "0010"; d2 <= "0101"; d3 <= "1001"; d4 <= "0000"; -- 952
    when "0000001110111001" => d1 <= "0011"; d2 <= "0101"; d3 <= "1001"; d4 <= "0000"; -- 953
    when "0000001110111010" => d1 <= "0100"; d2 <= "0101"; d3 <= "1001"; d4 <= "0000"; -- 954
    when "0000001110111011" => d1 <= "0101"; d2 <= "0101"; d3 <= "1001"; d4 <= "0000"; -- 955
    when "0000001110111100" => d1 <= "0110"; d2 <= "0101"; d3 <= "1001"; d4 <= "0000"; -- 956
    when "0000001110111101" => d1 <= "0111"; d2 <= "0101"; d3 <= "1001"; d4 <= "0000"; -- 957
    when "0000001110111110" => d1 <= "1000"; d2 <= "0101"; d3 <= "1001"; d4 <= "0000"; -- 958
    when "0000001110111111" => d1 <= "1001"; d2 <= "0101"; d3 <= "1001"; d4 <= "0000"; -- 959
    when "0000001111000000" => d1 <= "0000"; d2 <= "0110"; d3 <= "1001"; d4 <= "0000"; -- 960
    when "0000001111000001" => d1 <= "0001"; d2 <= "0110"; d3 <= "1001"; d4 <= "0000"; -- 961
    when "0000001111000010" => d1 <= "0010"; d2 <= "0110"; d3 <= "1001"; d4 <= "0000"; -- 962
    when "0000001111000011" => d1 <= "0011"; d2 <= "0110"; d3 <= "1001"; d4 <= "0000"; -- 963
    when "0000001111000100" => d1 <= "0100"; d2 <= "0110"; d3 <= "1001"; d4 <= "0000"; -- 964
    when "0000001111000101" => d1 <= "0101"; d2 <= "0110"; d3 <= "1001"; d4 <= "0000"; -- 965
    when "0000001111000110" => d1 <= "0110"; d2 <= "0110"; d3 <= "1001"; d4 <= "0000"; -- 966
    when "0000001111000111" => d1 <= "0111"; d2 <= "0110"; d3 <= "1001"; d4 <= "0000"; -- 967
    when "0000001111001000" => d1 <= "1000"; d2 <= "0110"; d3 <= "1001"; d4 <= "0000"; -- 968
    when "0000001111001001" => d1 <= "1001"; d2 <= "0110"; d3 <= "1001"; d4 <= "0000"; -- 969
    when "0000001111001010" => d1 <= "0000"; d2 <= "0111"; d3 <= "1001"; d4 <= "0000"; -- 970
    when "0000001111001011" => d1 <= "0001"; d2 <= "0111"; d3 <= "1001"; d4 <= "0000"; -- 971
    when "0000001111001100" => d1 <= "0010"; d2 <= "0111"; d3 <= "1001"; d4 <= "0000"; -- 972
    when "0000001111001101" => d1 <= "0011"; d2 <= "0111"; d3 <= "1001"; d4 <= "0000"; -- 973
    when "0000001111001110" => d1 <= "0100"; d2 <= "0111"; d3 <= "1001"; d4 <= "0000"; -- 974
    when "0000001111001111" => d1 <= "0101"; d2 <= "0111"; d3 <= "1001"; d4 <= "0000"; -- 975
    when "0000001111010000" => d1 <= "0110"; d2 <= "0111"; d3 <= "1001"; d4 <= "0000"; -- 976
    when "0000001111010001" => d1 <= "0111"; d2 <= "0111"; d3 <= "1001"; d4 <= "0000"; -- 977
    when "0000001111010010" => d1 <= "1000"; d2 <= "0111"; d3 <= "1001"; d4 <= "0000"; -- 978
    when "0000001111010011" => d1 <= "1001"; d2 <= "0111"; d3 <= "1001"; d4 <= "0000"; -- 979
    when "0000001111010100" => d1 <= "0000"; d2 <= "1000"; d3 <= "1001"; d4 <= "0000"; -- 980
    when "0000001111010101" => d1 <= "0001"; d2 <= "1000"; d3 <= "1001"; d4 <= "0000"; -- 981
    when "0000001111010110" => d1 <= "0010"; d2 <= "1000"; d3 <= "1001"; d4 <= "0000"; -- 982
    when "0000001111010111" => d1 <= "0011"; d2 <= "1000"; d3 <= "1001"; d4 <= "0000"; -- 983
    when "0000001111011000" => d1 <= "0100"; d2 <= "1000"; d3 <= "1001"; d4 <= "0000"; -- 984
    when "0000001111011001" => d1 <= "0101"; d2 <= "1000"; d3 <= "1001"; d4 <= "0000"; -- 985
    when "0000001111011010" => d1 <= "0110"; d2 <= "1000"; d3 <= "1001"; d4 <= "0000"; -- 986
    when "0000001111011011" => d1 <= "0111"; d2 <= "1000"; d3 <= "1001"; d4 <= "0000"; -- 987
    when "0000001111011100" => d1 <= "1000"; d2 <= "1000"; d3 <= "1001"; d4 <= "0000"; -- 988
    when "0000001111011101" => d1 <= "1001"; d2 <= "1000"; d3 <= "1001"; d4 <= "0000"; -- 989
    when "0000001111011110" => d1 <= "0000"; d2 <= "1001"; d3 <= "1001"; d4 <= "0000"; -- 990
    when "0000001111011111" => d1 <= "0001"; d2 <= "1001"; d3 <= "1001"; d4 <= "0000"; -- 991
    when "0000001111100000" => d1 <= "0010"; d2 <= "1001"; d3 <= "1001"; d4 <= "0000"; -- 992
    when "0000001111100001" => d1 <= "0011"; d2 <= "1001"; d3 <= "1001"; d4 <= "0000"; -- 993
    when "0000001111100010" => d1 <= "0100"; d2 <= "1001"; d3 <= "1001"; d4 <= "0000"; -- 994
    when "0000001111100011" => d1 <= "0101"; d2 <= "1001"; d3 <= "1001"; d4 <= "0000"; -- 995
    when "0000001111100100" => d1 <= "0110"; d2 <= "1001"; d3 <= "1001"; d4 <= "0000"; -- 996
    when "0000001111100101" => d1 <= "0111"; d2 <= "1001"; d3 <= "1001"; d4 <= "0000"; -- 997
    when "0000001111100110" => d1 <= "1000"; d2 <= "1001"; d3 <= "1001"; d4 <= "0000"; -- 998
    when "0000001111100111" => d1 <= "1001"; d2 <= "1001"; d3 <= "1001"; d4 <= "0000"; -- 999
    when "0000001111101000" => d1 <= "0000"; d2 <= "0000"; d3 <= "0000"; d4 <= "0001"; -- 1000
    when "0000001111101001" => d1 <= "0001"; d2 <= "0000"; d3 <= "0000"; d4 <= "0001"; -- 1001
    when "0000001111101010" => d1 <= "0010"; d2 <= "0000"; d3 <= "0000"; d4 <= "0001"; -- 1002
    when "0000001111101011" => d1 <= "0011"; d2 <= "0000"; d3 <= "0000"; d4 <= "0001"; -- 1003
    when "0000001111101100" => d1 <= "0100"; d2 <= "0000"; d3 <= "0000"; d4 <= "0001"; -- 1004
    when "0000001111101101" => d1 <= "0101"; d2 <= "0000"; d3 <= "0000"; d4 <= "0001"; -- 1005
    when "0000001111101110" => d1 <= "0110"; d2 <= "0000"; d3 <= "0000"; d4 <= "0001"; -- 1006
    when "0000001111101111" => d1 <= "0111"; d2 <= "0000"; d3 <= "0000"; d4 <= "0001"; -- 1007
    when "0000001111110000" => d1 <= "1000"; d2 <= "0000"; d3 <= "0000"; d4 <= "0001"; -- 1008
    when "0000001111110001" => d1 <= "1001"; d2 <= "0000"; d3 <= "0000"; d4 <= "0001"; -- 1009
    when "0000001111110010" => d1 <= "0000"; d2 <= "0001"; d3 <= "0000"; d4 <= "0001"; -- 1010
    when "0000001111110011" => d1 <= "0001"; d2 <= "0001"; d3 <= "0000"; d4 <= "0001"; -- 1011
    when "0000001111110100" => d1 <= "0010"; d2 <= "0001"; d3 <= "0000"; d4 <= "0001"; -- 1012
    when "0000001111110101" => d1 <= "0011"; d2 <= "0001"; d3 <= "0000"; d4 <= "0001"; -- 1013
    when "0000001111110110" => d1 <= "0100"; d2 <= "0001"; d3 <= "0000"; d4 <= "0001"; -- 1014
    when "0000001111110111" => d1 <= "0101"; d2 <= "0001"; d3 <= "0000"; d4 <= "0001"; -- 1015
    when "0000001111111000" => d1 <= "0110"; d2 <= "0001"; d3 <= "0000"; d4 <= "0001"; -- 1016
    when "0000001111111001" => d1 <= "0111"; d2 <= "0001"; d3 <= "0000"; d4 <= "0001"; -- 1017
    when "0000001111111010" => d1 <= "1000"; d2 <= "0001"; d3 <= "0000"; d4 <= "0001"; -- 1018
    when "0000001111111011" => d1 <= "1001"; d2 <= "0001"; d3 <= "0000"; d4 <= "0001"; -- 1019
    when "0000001111111100" => d1 <= "0000"; d2 <= "0010"; d3 <= "0000"; d4 <= "0001"; -- 1020
    when "0000001111111101" => d1 <= "0001"; d2 <= "0010"; d3 <= "0000"; d4 <= "0001"; -- 1021
    when "0000001111111110" => d1 <= "0010"; d2 <= "0010"; d3 <= "0000"; d4 <= "0001"; -- 1022
    when "0000001111111111" => d1 <= "0011"; d2 <= "0010"; d3 <= "0000"; d4 <= "0001"; -- 1023
    when "0000010000000000" => d1 <= "0100"; d2 <= "0010"; d3 <= "0000"; d4 <= "0001"; -- 1024
    when "0000010000000001" => d1 <= "0101"; d2 <= "0010"; d3 <= "0000"; d4 <= "0001"; -- 1025
    when "0000010000000010" => d1 <= "0110"; d2 <= "0010"; d3 <= "0000"; d4 <= "0001"; -- 1026
    when "0000010000000011" => d1 <= "0111"; d2 <= "0010"; d3 <= "0000"; d4 <= "0001"; -- 1027
    when "0000010000000100" => d1 <= "1000"; d2 <= "0010"; d3 <= "0000"; d4 <= "0001"; -- 1028
    when "0000010000000101" => d1 <= "1001"; d2 <= "0010"; d3 <= "0000"; d4 <= "0001"; -- 1029
    when "0000010000000110" => d1 <= "0000"; d2 <= "0011"; d3 <= "0000"; d4 <= "0001"; -- 1030
    when "0000010000000111" => d1 <= "0001"; d2 <= "0011"; d3 <= "0000"; d4 <= "0001"; -- 1031
    when "0000010000001000" => d1 <= "0010"; d2 <= "0011"; d3 <= "0000"; d4 <= "0001"; -- 1032
    when "0000010000001001" => d1 <= "0011"; d2 <= "0011"; d3 <= "0000"; d4 <= "0001"; -- 1033
    when "0000010000001010" => d1 <= "0100"; d2 <= "0011"; d3 <= "0000"; d4 <= "0001"; -- 1034
    when "0000010000001011" => d1 <= "0101"; d2 <= "0011"; d3 <= "0000"; d4 <= "0001"; -- 1035
    when "0000010000001100" => d1 <= "0110"; d2 <= "0011"; d3 <= "0000"; d4 <= "0001"; -- 1036
    when "0000010000001101" => d1 <= "0111"; d2 <= "0011"; d3 <= "0000"; d4 <= "0001"; -- 1037
    when "0000010000001110" => d1 <= "1000"; d2 <= "0011"; d3 <= "0000"; d4 <= "0001"; -- 1038
    when "0000010000001111" => d1 <= "1001"; d2 <= "0011"; d3 <= "0000"; d4 <= "0001"; -- 1039
    when "0000010000010000" => d1 <= "0000"; d2 <= "0100"; d3 <= "0000"; d4 <= "0001"; -- 1040
    when "0000010000010001" => d1 <= "0001"; d2 <= "0100"; d3 <= "0000"; d4 <= "0001"; -- 1041
    when "0000010000010010" => d1 <= "0010"; d2 <= "0100"; d3 <= "0000"; d4 <= "0001"; -- 1042
    when "0000010000010011" => d1 <= "0011"; d2 <= "0100"; d3 <= "0000"; d4 <= "0001"; -- 1043
    when "0000010000010100" => d1 <= "0100"; d2 <= "0100"; d3 <= "0000"; d4 <= "0001"; -- 1044
    when "0000010000010101" => d1 <= "0101"; d2 <= "0100"; d3 <= "0000"; d4 <= "0001"; -- 1045
    when "0000010000010110" => d1 <= "0110"; d2 <= "0100"; d3 <= "0000"; d4 <= "0001"; -- 1046
    when "0000010000010111" => d1 <= "0111"; d2 <= "0100"; d3 <= "0000"; d4 <= "0001"; -- 1047
    when "0000010000011000" => d1 <= "1000"; d2 <= "0100"; d3 <= "0000"; d4 <= "0001"; -- 1048
    when "0000010000011001" => d1 <= "1001"; d2 <= "0100"; d3 <= "0000"; d4 <= "0001"; -- 1049
    when "0000010000011010" => d1 <= "0000"; d2 <= "0101"; d3 <= "0000"; d4 <= "0001"; -- 1050
    when "0000010000011011" => d1 <= "0001"; d2 <= "0101"; d3 <= "0000"; d4 <= "0001"; -- 1051
    when "0000010000011100" => d1 <= "0010"; d2 <= "0101"; d3 <= "0000"; d4 <= "0001"; -- 1052
    when "0000010000011101" => d1 <= "0011"; d2 <= "0101"; d3 <= "0000"; d4 <= "0001"; -- 1053
    when "0000010000011110" => d1 <= "0100"; d2 <= "0101"; d3 <= "0000"; d4 <= "0001"; -- 1054
    when "0000010000011111" => d1 <= "0101"; d2 <= "0101"; d3 <= "0000"; d4 <= "0001"; -- 1055
    when "0000010000100000" => d1 <= "0110"; d2 <= "0101"; d3 <= "0000"; d4 <= "0001"; -- 1056
    when "0000010000100001" => d1 <= "0111"; d2 <= "0101"; d3 <= "0000"; d4 <= "0001"; -- 1057
    when "0000010000100010" => d1 <= "1000"; d2 <= "0101"; d3 <= "0000"; d4 <= "0001"; -- 1058
    when "0000010000100011" => d1 <= "1001"; d2 <= "0101"; d3 <= "0000"; d4 <= "0001"; -- 1059
    when "0000010000100100" => d1 <= "0000"; d2 <= "0110"; d3 <= "0000"; d4 <= "0001"; -- 1060
    when "0000010000100101" => d1 <= "0001"; d2 <= "0110"; d3 <= "0000"; d4 <= "0001"; -- 1061
    when "0000010000100110" => d1 <= "0010"; d2 <= "0110"; d3 <= "0000"; d4 <= "0001"; -- 1062
    when "0000010000100111" => d1 <= "0011"; d2 <= "0110"; d3 <= "0000"; d4 <= "0001"; -- 1063
    when "0000010000101000" => d1 <= "0100"; d2 <= "0110"; d3 <= "0000"; d4 <= "0001"; -- 1064
    when "0000010000101001" => d1 <= "0101"; d2 <= "0110"; d3 <= "0000"; d4 <= "0001"; -- 1065
    when "0000010000101010" => d1 <= "0110"; d2 <= "0110"; d3 <= "0000"; d4 <= "0001"; -- 1066
    when "0000010000101011" => d1 <= "0111"; d2 <= "0110"; d3 <= "0000"; d4 <= "0001"; -- 1067
    when "0000010000101100" => d1 <= "1000"; d2 <= "0110"; d3 <= "0000"; d4 <= "0001"; -- 1068
    when "0000010000101101" => d1 <= "1001"; d2 <= "0110"; d3 <= "0000"; d4 <= "0001"; -- 1069
    when "0000010000101110" => d1 <= "0000"; d2 <= "0111"; d3 <= "0000"; d4 <= "0001"; -- 1070
    when "0000010000101111" => d1 <= "0001"; d2 <= "0111"; d3 <= "0000"; d4 <= "0001"; -- 1071
    when "0000010000110000" => d1 <= "0010"; d2 <= "0111"; d3 <= "0000"; d4 <= "0001"; -- 1072
    when "0000010000110001" => d1 <= "0011"; d2 <= "0111"; d3 <= "0000"; d4 <= "0001"; -- 1073
    when "0000010000110010" => d1 <= "0100"; d2 <= "0111"; d3 <= "0000"; d4 <= "0001"; -- 1074
    when "0000010000110011" => d1 <= "0101"; d2 <= "0111"; d3 <= "0000"; d4 <= "0001"; -- 1075
    when "0000010000110100" => d1 <= "0110"; d2 <= "0111"; d3 <= "0000"; d4 <= "0001"; -- 1076
    when "0000010000110101" => d1 <= "0111"; d2 <= "0111"; d3 <= "0000"; d4 <= "0001"; -- 1077
    when "0000010000110110" => d1 <= "1000"; d2 <= "0111"; d3 <= "0000"; d4 <= "0001"; -- 1078
    when "0000010000110111" => d1 <= "1001"; d2 <= "0111"; d3 <= "0000"; d4 <= "0001"; -- 1079
    when "0000010000111000" => d1 <= "0000"; d2 <= "1000"; d3 <= "0000"; d4 <= "0001"; -- 1080
    when "0000010000111001" => d1 <= "0001"; d2 <= "1000"; d3 <= "0000"; d4 <= "0001"; -- 1081
    when "0000010000111010" => d1 <= "0010"; d2 <= "1000"; d3 <= "0000"; d4 <= "0001"; -- 1082
    when "0000010000111011" => d1 <= "0011"; d2 <= "1000"; d3 <= "0000"; d4 <= "0001"; -- 1083
    when "0000010000111100" => d1 <= "0100"; d2 <= "1000"; d3 <= "0000"; d4 <= "0001"; -- 1084
    when "0000010000111101" => d1 <= "0101"; d2 <= "1000"; d3 <= "0000"; d4 <= "0001"; -- 1085
    when "0000010000111110" => d1 <= "0110"; d2 <= "1000"; d3 <= "0000"; d4 <= "0001"; -- 1086
    when "0000010000111111" => d1 <= "0111"; d2 <= "1000"; d3 <= "0000"; d4 <= "0001"; -- 1087
    when "0000010001000000" => d1 <= "1000"; d2 <= "1000"; d3 <= "0000"; d4 <= "0001"; -- 1088
    when "0000010001000001" => d1 <= "1001"; d2 <= "1000"; d3 <= "0000"; d4 <= "0001"; -- 1089
    when "0000010001000010" => d1 <= "0000"; d2 <= "1001"; d3 <= "0000"; d4 <= "0001"; -- 1090
    when "0000010001000011" => d1 <= "0001"; d2 <= "1001"; d3 <= "0000"; d4 <= "0001"; -- 1091
    when "0000010001000100" => d1 <= "0010"; d2 <= "1001"; d3 <= "0000"; d4 <= "0001"; -- 1092
    when "0000010001000101" => d1 <= "0011"; d2 <= "1001"; d3 <= "0000"; d4 <= "0001"; -- 1093
    when "0000010001000110" => d1 <= "0100"; d2 <= "1001"; d3 <= "0000"; d4 <= "0001"; -- 1094
    when "0000010001000111" => d1 <= "0101"; d2 <= "1001"; d3 <= "0000"; d4 <= "0001"; -- 1095
    when "0000010001001000" => d1 <= "0110"; d2 <= "1001"; d3 <= "0000"; d4 <= "0001"; -- 1096
    when "0000010001001001" => d1 <= "0111"; d2 <= "1001"; d3 <= "0000"; d4 <= "0001"; -- 1097
    when "0000010001001010" => d1 <= "1000"; d2 <= "1001"; d3 <= "0000"; d4 <= "0001"; -- 1098
    when "0000010001001011" => d1 <= "1001"; d2 <= "1001"; d3 <= "0000"; d4 <= "0001"; -- 1099
    when "0000010001001100" => d1 <= "0000"; d2 <= "0000"; d3 <= "0001"; d4 <= "0001"; -- 1100
    when "0000010001001101" => d1 <= "0001"; d2 <= "0000"; d3 <= "0001"; d4 <= "0001"; -- 1101
    when "0000010001001110" => d1 <= "0010"; d2 <= "0000"; d3 <= "0001"; d4 <= "0001"; -- 1102
    when "0000010001001111" => d1 <= "0011"; d2 <= "0000"; d3 <= "0001"; d4 <= "0001"; -- 1103
    when "0000010001010000" => d1 <= "0100"; d2 <= "0000"; d3 <= "0001"; d4 <= "0001"; -- 1104
    when "0000010001010001" => d1 <= "0101"; d2 <= "0000"; d3 <= "0001"; d4 <= "0001"; -- 1105
    when "0000010001010010" => d1 <= "0110"; d2 <= "0000"; d3 <= "0001"; d4 <= "0001"; -- 1106
    when "0000010001010011" => d1 <= "0111"; d2 <= "0000"; d3 <= "0001"; d4 <= "0001"; -- 1107
    when "0000010001010100" => d1 <= "1000"; d2 <= "0000"; d3 <= "0001"; d4 <= "0001"; -- 1108
    when "0000010001010101" => d1 <= "1001"; d2 <= "0000"; d3 <= "0001"; d4 <= "0001"; -- 1109
    when "0000010001010110" => d1 <= "0000"; d2 <= "0001"; d3 <= "0001"; d4 <= "0001"; -- 1110
    when "0000010001010111" => d1 <= "0001"; d2 <= "0001"; d3 <= "0001"; d4 <= "0001"; -- 1111
    when "0000010001011000" => d1 <= "0010"; d2 <= "0001"; d3 <= "0001"; d4 <= "0001"; -- 1112
    when "0000010001011001" => d1 <= "0011"; d2 <= "0001"; d3 <= "0001"; d4 <= "0001"; -- 1113
    when "0000010001011010" => d1 <= "0100"; d2 <= "0001"; d3 <= "0001"; d4 <= "0001"; -- 1114
    when "0000010001011011" => d1 <= "0101"; d2 <= "0001"; d3 <= "0001"; d4 <= "0001"; -- 1115
    when "0000010001011100" => d1 <= "0110"; d2 <= "0001"; d3 <= "0001"; d4 <= "0001"; -- 1116
    when "0000010001011101" => d1 <= "0111"; d2 <= "0001"; d3 <= "0001"; d4 <= "0001"; -- 1117
    when "0000010001011110" => d1 <= "1000"; d2 <= "0001"; d3 <= "0001"; d4 <= "0001"; -- 1118
    when "0000010001011111" => d1 <= "1001"; d2 <= "0001"; d3 <= "0001"; d4 <= "0001"; -- 1119
    when "0000010001100000" => d1 <= "0000"; d2 <= "0010"; d3 <= "0001"; d4 <= "0001"; -- 1120
    when "0000010001100001" => d1 <= "0001"; d2 <= "0010"; d3 <= "0001"; d4 <= "0001"; -- 1121
    when "0000010001100010" => d1 <= "0010"; d2 <= "0010"; d3 <= "0001"; d4 <= "0001"; -- 1122
    when "0000010001100011" => d1 <= "0011"; d2 <= "0010"; d3 <= "0001"; d4 <= "0001"; -- 1123
    when "0000010001100100" => d1 <= "0100"; d2 <= "0010"; d3 <= "0001"; d4 <= "0001"; -- 1124
    when "0000010001100101" => d1 <= "0101"; d2 <= "0010"; d3 <= "0001"; d4 <= "0001"; -- 1125
    when "0000010001100110" => d1 <= "0110"; d2 <= "0010"; d3 <= "0001"; d4 <= "0001"; -- 1126
    when "0000010001100111" => d1 <= "0111"; d2 <= "0010"; d3 <= "0001"; d4 <= "0001"; -- 1127
    when "0000010001101000" => d1 <= "1000"; d2 <= "0010"; d3 <= "0001"; d4 <= "0001"; -- 1128
    when "0000010001101001" => d1 <= "1001"; d2 <= "0010"; d3 <= "0001"; d4 <= "0001"; -- 1129
    when "0000010001101010" => d1 <= "0000"; d2 <= "0011"; d3 <= "0001"; d4 <= "0001"; -- 1130
    when "0000010001101011" => d1 <= "0001"; d2 <= "0011"; d3 <= "0001"; d4 <= "0001"; -- 1131
    when "0000010001101100" => d1 <= "0010"; d2 <= "0011"; d3 <= "0001"; d4 <= "0001"; -- 1132
    when "0000010001101101" => d1 <= "0011"; d2 <= "0011"; d3 <= "0001"; d4 <= "0001"; -- 1133
    when "0000010001101110" => d1 <= "0100"; d2 <= "0011"; d3 <= "0001"; d4 <= "0001"; -- 1134
    when "0000010001101111" => d1 <= "0101"; d2 <= "0011"; d3 <= "0001"; d4 <= "0001"; -- 1135
    when "0000010001110000" => d1 <= "0110"; d2 <= "0011"; d3 <= "0001"; d4 <= "0001"; -- 1136
    when "0000010001110001" => d1 <= "0111"; d2 <= "0011"; d3 <= "0001"; d4 <= "0001"; -- 1137
    when "0000010001110010" => d1 <= "1000"; d2 <= "0011"; d3 <= "0001"; d4 <= "0001"; -- 1138
    when "0000010001110011" => d1 <= "1001"; d2 <= "0011"; d3 <= "0001"; d4 <= "0001"; -- 1139
    when "0000010001110100" => d1 <= "0000"; d2 <= "0100"; d3 <= "0001"; d4 <= "0001"; -- 1140
    when "0000010001110101" => d1 <= "0001"; d2 <= "0100"; d3 <= "0001"; d4 <= "0001"; -- 1141
    when "0000010001110110" => d1 <= "0010"; d2 <= "0100"; d3 <= "0001"; d4 <= "0001"; -- 1142
    when "0000010001110111" => d1 <= "0011"; d2 <= "0100"; d3 <= "0001"; d4 <= "0001"; -- 1143
    when "0000010001111000" => d1 <= "0100"; d2 <= "0100"; d3 <= "0001"; d4 <= "0001"; -- 1144
    when "0000010001111001" => d1 <= "0101"; d2 <= "0100"; d3 <= "0001"; d4 <= "0001"; -- 1145
    when "0000010001111010" => d1 <= "0110"; d2 <= "0100"; d3 <= "0001"; d4 <= "0001"; -- 1146
    when "0000010001111011" => d1 <= "0111"; d2 <= "0100"; d3 <= "0001"; d4 <= "0001"; -- 1147
    when "0000010001111100" => d1 <= "1000"; d2 <= "0100"; d3 <= "0001"; d4 <= "0001"; -- 1148
    when "0000010001111101" => d1 <= "1001"; d2 <= "0100"; d3 <= "0001"; d4 <= "0001"; -- 1149
    when "0000010001111110" => d1 <= "0000"; d2 <= "0101"; d3 <= "0001"; d4 <= "0001"; -- 1150
    when "0000010001111111" => d1 <= "0001"; d2 <= "0101"; d3 <= "0001"; d4 <= "0001"; -- 1151
    when "0000010010000000" => d1 <= "0010"; d2 <= "0101"; d3 <= "0001"; d4 <= "0001"; -- 1152
    when "0000010010000001" => d1 <= "0011"; d2 <= "0101"; d3 <= "0001"; d4 <= "0001"; -- 1153
    when "0000010010000010" => d1 <= "0100"; d2 <= "0101"; d3 <= "0001"; d4 <= "0001"; -- 1154
    when "0000010010000011" => d1 <= "0101"; d2 <= "0101"; d3 <= "0001"; d4 <= "0001"; -- 1155
    when "0000010010000100" => d1 <= "0110"; d2 <= "0101"; d3 <= "0001"; d4 <= "0001"; -- 1156
    when "0000010010000101" => d1 <= "0111"; d2 <= "0101"; d3 <= "0001"; d4 <= "0001"; -- 1157
    when "0000010010000110" => d1 <= "1000"; d2 <= "0101"; d3 <= "0001"; d4 <= "0001"; -- 1158
    when "0000010010000111" => d1 <= "1001"; d2 <= "0101"; d3 <= "0001"; d4 <= "0001"; -- 1159
    when "0000010010001000" => d1 <= "0000"; d2 <= "0110"; d3 <= "0001"; d4 <= "0001"; -- 1160
    when "0000010010001001" => d1 <= "0001"; d2 <= "0110"; d3 <= "0001"; d4 <= "0001"; -- 1161
    when "0000010010001010" => d1 <= "0010"; d2 <= "0110"; d3 <= "0001"; d4 <= "0001"; -- 1162
    when "0000010010001011" => d1 <= "0011"; d2 <= "0110"; d3 <= "0001"; d4 <= "0001"; -- 1163
    when "0000010010001100" => d1 <= "0100"; d2 <= "0110"; d3 <= "0001"; d4 <= "0001"; -- 1164
    when "0000010010001101" => d1 <= "0101"; d2 <= "0110"; d3 <= "0001"; d4 <= "0001"; -- 1165
    when "0000010010001110" => d1 <= "0110"; d2 <= "0110"; d3 <= "0001"; d4 <= "0001"; -- 1166
    when "0000010010001111" => d1 <= "0111"; d2 <= "0110"; d3 <= "0001"; d4 <= "0001"; -- 1167
    when "0000010010010000" => d1 <= "1000"; d2 <= "0110"; d3 <= "0001"; d4 <= "0001"; -- 1168
    when "0000010010010001" => d1 <= "1001"; d2 <= "0110"; d3 <= "0001"; d4 <= "0001"; -- 1169
    when "0000010010010010" => d1 <= "0000"; d2 <= "0111"; d3 <= "0001"; d4 <= "0001"; -- 1170
    when "0000010010010011" => d1 <= "0001"; d2 <= "0111"; d3 <= "0001"; d4 <= "0001"; -- 1171
    when "0000010010010100" => d1 <= "0010"; d2 <= "0111"; d3 <= "0001"; d4 <= "0001"; -- 1172
    when "0000010010010101" => d1 <= "0011"; d2 <= "0111"; d3 <= "0001"; d4 <= "0001"; -- 1173
    when "0000010010010110" => d1 <= "0100"; d2 <= "0111"; d3 <= "0001"; d4 <= "0001"; -- 1174
    when "0000010010010111" => d1 <= "0101"; d2 <= "0111"; d3 <= "0001"; d4 <= "0001"; -- 1175
    when "0000010010011000" => d1 <= "0110"; d2 <= "0111"; d3 <= "0001"; d4 <= "0001"; -- 1176
    when "0000010010011001" => d1 <= "0111"; d2 <= "0111"; d3 <= "0001"; d4 <= "0001"; -- 1177
    when "0000010010011010" => d1 <= "1000"; d2 <= "0111"; d3 <= "0001"; d4 <= "0001"; -- 1178
    when "0000010010011011" => d1 <= "1001"; d2 <= "0111"; d3 <= "0001"; d4 <= "0001"; -- 1179
    when "0000010010011100" => d1 <= "0000"; d2 <= "1000"; d3 <= "0001"; d4 <= "0001"; -- 1180
    when "0000010010011101" => d1 <= "0001"; d2 <= "1000"; d3 <= "0001"; d4 <= "0001"; -- 1181
    when "0000010010011110" => d1 <= "0010"; d2 <= "1000"; d3 <= "0001"; d4 <= "0001"; -- 1182
    when "0000010010011111" => d1 <= "0011"; d2 <= "1000"; d3 <= "0001"; d4 <= "0001"; -- 1183
    when "0000010010100000" => d1 <= "0100"; d2 <= "1000"; d3 <= "0001"; d4 <= "0001"; -- 1184
    when "0000010010100001" => d1 <= "0101"; d2 <= "1000"; d3 <= "0001"; d4 <= "0001"; -- 1185
    when "0000010010100010" => d1 <= "0110"; d2 <= "1000"; d3 <= "0001"; d4 <= "0001"; -- 1186
    when "0000010010100011" => d1 <= "0111"; d2 <= "1000"; d3 <= "0001"; d4 <= "0001"; -- 1187
    when "0000010010100100" => d1 <= "1000"; d2 <= "1000"; d3 <= "0001"; d4 <= "0001"; -- 1188
    when "0000010010100101" => d1 <= "1001"; d2 <= "1000"; d3 <= "0001"; d4 <= "0001"; -- 1189
    when "0000010010100110" => d1 <= "0000"; d2 <= "1001"; d3 <= "0001"; d4 <= "0001"; -- 1190
    when "0000010010100111" => d1 <= "0001"; d2 <= "1001"; d3 <= "0001"; d4 <= "0001"; -- 1191
    when "0000010010101000" => d1 <= "0010"; d2 <= "1001"; d3 <= "0001"; d4 <= "0001"; -- 1192
    when "0000010010101001" => d1 <= "0011"; d2 <= "1001"; d3 <= "0001"; d4 <= "0001"; -- 1193
    when "0000010010101010" => d1 <= "0100"; d2 <= "1001"; d3 <= "0001"; d4 <= "0001"; -- 1194
    when "0000010010101011" => d1 <= "0101"; d2 <= "1001"; d3 <= "0001"; d4 <= "0001"; -- 1195
    when "0000010010101100" => d1 <= "0110"; d2 <= "1001"; d3 <= "0001"; d4 <= "0001"; -- 1196
    when "0000010010101101" => d1 <= "0111"; d2 <= "1001"; d3 <= "0001"; d4 <= "0001"; -- 1197
    when "0000010010101110" => d1 <= "1000"; d2 <= "1001"; d3 <= "0001"; d4 <= "0001"; -- 1198
    when "0000010010101111" => d1 <= "1001"; d2 <= "1001"; d3 <= "0001"; d4 <= "0001"; -- 1199
    when "0000010010110000" => d1 <= "0000"; d2 <= "0000"; d3 <= "0010"; d4 <= "0001"; -- 1200
    when "0000010010110001" => d1 <= "0001"; d2 <= "0000"; d3 <= "0010"; d4 <= "0001"; -- 1201
    when "0000010010110010" => d1 <= "0010"; d2 <= "0000"; d3 <= "0010"; d4 <= "0001"; -- 1202
    when "0000010010110011" => d1 <= "0011"; d2 <= "0000"; d3 <= "0010"; d4 <= "0001"; -- 1203
    when "0000010010110100" => d1 <= "0100"; d2 <= "0000"; d3 <= "0010"; d4 <= "0001"; -- 1204
    when "0000010010110101" => d1 <= "0101"; d2 <= "0000"; d3 <= "0010"; d4 <= "0001"; -- 1205
    when "0000010010110110" => d1 <= "0110"; d2 <= "0000"; d3 <= "0010"; d4 <= "0001"; -- 1206
    when "0000010010110111" => d1 <= "0111"; d2 <= "0000"; d3 <= "0010"; d4 <= "0001"; -- 1207
    when "0000010010111000" => d1 <= "1000"; d2 <= "0000"; d3 <= "0010"; d4 <= "0001"; -- 1208
    when "0000010010111001" => d1 <= "1001"; d2 <= "0000"; d3 <= "0010"; d4 <= "0001"; -- 1209
    when "0000010010111010" => d1 <= "0000"; d2 <= "0001"; d3 <= "0010"; d4 <= "0001"; -- 1210
    when "0000010010111011" => d1 <= "0001"; d2 <= "0001"; d3 <= "0010"; d4 <= "0001"; -- 1211
    when "0000010010111100" => d1 <= "0010"; d2 <= "0001"; d3 <= "0010"; d4 <= "0001"; -- 1212
    when "0000010010111101" => d1 <= "0011"; d2 <= "0001"; d3 <= "0010"; d4 <= "0001"; -- 1213
    when "0000010010111110" => d1 <= "0100"; d2 <= "0001"; d3 <= "0010"; d4 <= "0001"; -- 1214
    when "0000010010111111" => d1 <= "0101"; d2 <= "0001"; d3 <= "0010"; d4 <= "0001"; -- 1215
    when "0000010011000000" => d1 <= "0110"; d2 <= "0001"; d3 <= "0010"; d4 <= "0001"; -- 1216
    when "0000010011000001" => d1 <= "0111"; d2 <= "0001"; d3 <= "0010"; d4 <= "0001"; -- 1217
    when "0000010011000010" => d1 <= "1000"; d2 <= "0001"; d3 <= "0010"; d4 <= "0001"; -- 1218
    when "0000010011000011" => d1 <= "1001"; d2 <= "0001"; d3 <= "0010"; d4 <= "0001"; -- 1219
    when "0000010011000100" => d1 <= "0000"; d2 <= "0010"; d3 <= "0010"; d4 <= "0001"; -- 1220
    when "0000010011000101" => d1 <= "0001"; d2 <= "0010"; d3 <= "0010"; d4 <= "0001"; -- 1221
    when "0000010011000110" => d1 <= "0010"; d2 <= "0010"; d3 <= "0010"; d4 <= "0001"; -- 1222
    when "0000010011000111" => d1 <= "0011"; d2 <= "0010"; d3 <= "0010"; d4 <= "0001"; -- 1223
    when "0000010011001000" => d1 <= "0100"; d2 <= "0010"; d3 <= "0010"; d4 <= "0001"; -- 1224
    when "0000010011001001" => d1 <= "0101"; d2 <= "0010"; d3 <= "0010"; d4 <= "0001"; -- 1225
    when "0000010011001010" => d1 <= "0110"; d2 <= "0010"; d3 <= "0010"; d4 <= "0001"; -- 1226
    when "0000010011001011" => d1 <= "0111"; d2 <= "0010"; d3 <= "0010"; d4 <= "0001"; -- 1227
    when "0000010011001100" => d1 <= "1000"; d2 <= "0010"; d3 <= "0010"; d4 <= "0001"; -- 1228
    when "0000010011001101" => d1 <= "1001"; d2 <= "0010"; d3 <= "0010"; d4 <= "0001"; -- 1229
    when "0000010011001110" => d1 <= "0000"; d2 <= "0011"; d3 <= "0010"; d4 <= "0001"; -- 1230
    when "0000010011001111" => d1 <= "0001"; d2 <= "0011"; d3 <= "0010"; d4 <= "0001"; -- 1231
    when "0000010011010000" => d1 <= "0010"; d2 <= "0011"; d3 <= "0010"; d4 <= "0001"; -- 1232
    when "0000010011010001" => d1 <= "0011"; d2 <= "0011"; d3 <= "0010"; d4 <= "0001"; -- 1233
    when "0000010011010010" => d1 <= "0100"; d2 <= "0011"; d3 <= "0010"; d4 <= "0001"; -- 1234
    when "0000010011010011" => d1 <= "0101"; d2 <= "0011"; d3 <= "0010"; d4 <= "0001"; -- 1235
    when "0000010011010100" => d1 <= "0110"; d2 <= "0011"; d3 <= "0010"; d4 <= "0001"; -- 1236
    when "0000010011010101" => d1 <= "0111"; d2 <= "0011"; d3 <= "0010"; d4 <= "0001"; -- 1237
    when "0000010011010110" => d1 <= "1000"; d2 <= "0011"; d3 <= "0010"; d4 <= "0001"; -- 1238
    when "0000010011010111" => d1 <= "1001"; d2 <= "0011"; d3 <= "0010"; d4 <= "0001"; -- 1239
    when "0000010011011000" => d1 <= "0000"; d2 <= "0100"; d3 <= "0010"; d4 <= "0001"; -- 1240
    when "0000010011011001" => d1 <= "0001"; d2 <= "0100"; d3 <= "0010"; d4 <= "0001"; -- 1241
    when "0000010011011010" => d1 <= "0010"; d2 <= "0100"; d3 <= "0010"; d4 <= "0001"; -- 1242
    when "0000010011011011" => d1 <= "0011"; d2 <= "0100"; d3 <= "0010"; d4 <= "0001"; -- 1243
    when "0000010011011100" => d1 <= "0100"; d2 <= "0100"; d3 <= "0010"; d4 <= "0001"; -- 1244
    when "0000010011011101" => d1 <= "0101"; d2 <= "0100"; d3 <= "0010"; d4 <= "0001"; -- 1245
    when "0000010011011110" => d1 <= "0110"; d2 <= "0100"; d3 <= "0010"; d4 <= "0001"; -- 1246
    when "0000010011011111" => d1 <= "0111"; d2 <= "0100"; d3 <= "0010"; d4 <= "0001"; -- 1247
    when "0000010011100000" => d1 <= "1000"; d2 <= "0100"; d3 <= "0010"; d4 <= "0001"; -- 1248
    when "0000010011100001" => d1 <= "1001"; d2 <= "0100"; d3 <= "0010"; d4 <= "0001"; -- 1249
    when "0000010011100010" => d1 <= "0000"; d2 <= "0101"; d3 <= "0010"; d4 <= "0001"; -- 1250
    when "0000010011100011" => d1 <= "0001"; d2 <= "0101"; d3 <= "0010"; d4 <= "0001"; -- 1251
    when "0000010011100100" => d1 <= "0010"; d2 <= "0101"; d3 <= "0010"; d4 <= "0001"; -- 1252
    when "0000010011100101" => d1 <= "0011"; d2 <= "0101"; d3 <= "0010"; d4 <= "0001"; -- 1253
    when "0000010011100110" => d1 <= "0100"; d2 <= "0101"; d3 <= "0010"; d4 <= "0001"; -- 1254
    when "0000010011100111" => d1 <= "0101"; d2 <= "0101"; d3 <= "0010"; d4 <= "0001"; -- 1255
    when "0000010011101000" => d1 <= "0110"; d2 <= "0101"; d3 <= "0010"; d4 <= "0001"; -- 1256
    when "0000010011101001" => d1 <= "0111"; d2 <= "0101"; d3 <= "0010"; d4 <= "0001"; -- 1257
    when "0000010011101010" => d1 <= "1000"; d2 <= "0101"; d3 <= "0010"; d4 <= "0001"; -- 1258
    when "0000010011101011" => d1 <= "1001"; d2 <= "0101"; d3 <= "0010"; d4 <= "0001"; -- 1259
    when "0000010011101100" => d1 <= "0000"; d2 <= "0110"; d3 <= "0010"; d4 <= "0001"; -- 1260
    when "0000010011101101" => d1 <= "0001"; d2 <= "0110"; d3 <= "0010"; d4 <= "0001"; -- 1261
    when "0000010011101110" => d1 <= "0010"; d2 <= "0110"; d3 <= "0010"; d4 <= "0001"; -- 1262
    when "0000010011101111" => d1 <= "0011"; d2 <= "0110"; d3 <= "0010"; d4 <= "0001"; -- 1263
    when "0000010011110000" => d1 <= "0100"; d2 <= "0110"; d3 <= "0010"; d4 <= "0001"; -- 1264
    when "0000010011110001" => d1 <= "0101"; d2 <= "0110"; d3 <= "0010"; d4 <= "0001"; -- 1265
    when "0000010011110010" => d1 <= "0110"; d2 <= "0110"; d3 <= "0010"; d4 <= "0001"; -- 1266
    when "0000010011110011" => d1 <= "0111"; d2 <= "0110"; d3 <= "0010"; d4 <= "0001"; -- 1267
    when "0000010011110100" => d1 <= "1000"; d2 <= "0110"; d3 <= "0010"; d4 <= "0001"; -- 1268
    when "0000010011110101" => d1 <= "1001"; d2 <= "0110"; d3 <= "0010"; d4 <= "0001"; -- 1269
    when "0000010011110110" => d1 <= "0000"; d2 <= "0111"; d3 <= "0010"; d4 <= "0001"; -- 1270
    when "0000010011110111" => d1 <= "0001"; d2 <= "0111"; d3 <= "0010"; d4 <= "0001"; -- 1271
    when "0000010011111000" => d1 <= "0010"; d2 <= "0111"; d3 <= "0010"; d4 <= "0001"; -- 1272
    when "0000010011111001" => d1 <= "0011"; d2 <= "0111"; d3 <= "0010"; d4 <= "0001"; -- 1273
    when "0000010011111010" => d1 <= "0100"; d2 <= "0111"; d3 <= "0010"; d4 <= "0001"; -- 1274
    when "0000010011111011" => d1 <= "0101"; d2 <= "0111"; d3 <= "0010"; d4 <= "0001"; -- 1275
    when "0000010011111100" => d1 <= "0110"; d2 <= "0111"; d3 <= "0010"; d4 <= "0001"; -- 1276
    when "0000010011111101" => d1 <= "0111"; d2 <= "0111"; d3 <= "0010"; d4 <= "0001"; -- 1277
    when "0000010011111110" => d1 <= "1000"; d2 <= "0111"; d3 <= "0010"; d4 <= "0001"; -- 1278
    when "0000010011111111" => d1 <= "1001"; d2 <= "0111"; d3 <= "0010"; d4 <= "0001"; -- 1279
    when "0000010100000000" => d1 <= "0000"; d2 <= "1000"; d3 <= "0010"; d4 <= "0001"; -- 1280
    when "0000010100000001" => d1 <= "0001"; d2 <= "1000"; d3 <= "0010"; d4 <= "0001"; -- 1281
    when "0000010100000010" => d1 <= "0010"; d2 <= "1000"; d3 <= "0010"; d4 <= "0001"; -- 1282
    when "0000010100000011" => d1 <= "0011"; d2 <= "1000"; d3 <= "0010"; d4 <= "0001"; -- 1283
    when "0000010100000100" => d1 <= "0100"; d2 <= "1000"; d3 <= "0010"; d4 <= "0001"; -- 1284
    when "0000010100000101" => d1 <= "0101"; d2 <= "1000"; d3 <= "0010"; d4 <= "0001"; -- 1285
    when "0000010100000110" => d1 <= "0110"; d2 <= "1000"; d3 <= "0010"; d4 <= "0001"; -- 1286
    when "0000010100000111" => d1 <= "0111"; d2 <= "1000"; d3 <= "0010"; d4 <= "0001"; -- 1287
    when "0000010100001000" => d1 <= "1000"; d2 <= "1000"; d3 <= "0010"; d4 <= "0001"; -- 1288
    when "0000010100001001" => d1 <= "1001"; d2 <= "1000"; d3 <= "0010"; d4 <= "0001"; -- 1289
    when "0000010100001010" => d1 <= "0000"; d2 <= "1001"; d3 <= "0010"; d4 <= "0001"; -- 1290
    when "0000010100001011" => d1 <= "0001"; d2 <= "1001"; d3 <= "0010"; d4 <= "0001"; -- 1291
    when "0000010100001100" => d1 <= "0010"; d2 <= "1001"; d3 <= "0010"; d4 <= "0001"; -- 1292
    when "0000010100001101" => d1 <= "0011"; d2 <= "1001"; d3 <= "0010"; d4 <= "0001"; -- 1293
    when "0000010100001110" => d1 <= "0100"; d2 <= "1001"; d3 <= "0010"; d4 <= "0001"; -- 1294
    when "0000010100001111" => d1 <= "0101"; d2 <= "1001"; d3 <= "0010"; d4 <= "0001"; -- 1295
    when "0000010100010000" => d1 <= "0110"; d2 <= "1001"; d3 <= "0010"; d4 <= "0001"; -- 1296
    when "0000010100010001" => d1 <= "0111"; d2 <= "1001"; d3 <= "0010"; d4 <= "0001"; -- 1297
    when "0000010100010010" => d1 <= "1000"; d2 <= "1001"; d3 <= "0010"; d4 <= "0001"; -- 1298
    when "0000010100010011" => d1 <= "1001"; d2 <= "1001"; d3 <= "0010"; d4 <= "0001"; -- 1299
    when "0000010100010100" => d1 <= "0000"; d2 <= "0000"; d3 <= "0011"; d4 <= "0001"; -- 1300
    when "0000010100010101" => d1 <= "0001"; d2 <= "0000"; d3 <= "0011"; d4 <= "0001"; -- 1301
    when "0000010100010110" => d1 <= "0010"; d2 <= "0000"; d3 <= "0011"; d4 <= "0001"; -- 1302
    when "0000010100010111" => d1 <= "0011"; d2 <= "0000"; d3 <= "0011"; d4 <= "0001"; -- 1303
    when "0000010100011000" => d1 <= "0100"; d2 <= "0000"; d3 <= "0011"; d4 <= "0001"; -- 1304
    when "0000010100011001" => d1 <= "0101"; d2 <= "0000"; d3 <= "0011"; d4 <= "0001"; -- 1305
    when "0000010100011010" => d1 <= "0110"; d2 <= "0000"; d3 <= "0011"; d4 <= "0001"; -- 1306
    when "0000010100011011" => d1 <= "0111"; d2 <= "0000"; d3 <= "0011"; d4 <= "0001"; -- 1307
    when "0000010100011100" => d1 <= "1000"; d2 <= "0000"; d3 <= "0011"; d4 <= "0001"; -- 1308
    when "0000010100011101" => d1 <= "1001"; d2 <= "0000"; d3 <= "0011"; d4 <= "0001"; -- 1309
    when "0000010100011110" => d1 <= "0000"; d2 <= "0001"; d3 <= "0011"; d4 <= "0001"; -- 1310
    when "0000010100011111" => d1 <= "0001"; d2 <= "0001"; d3 <= "0011"; d4 <= "0001"; -- 1311
    when "0000010100100000" => d1 <= "0010"; d2 <= "0001"; d3 <= "0011"; d4 <= "0001"; -- 1312
    when "0000010100100001" => d1 <= "0011"; d2 <= "0001"; d3 <= "0011"; d4 <= "0001"; -- 1313
    when "0000010100100010" => d1 <= "0100"; d2 <= "0001"; d3 <= "0011"; d4 <= "0001"; -- 1314
    when "0000010100100011" => d1 <= "0101"; d2 <= "0001"; d3 <= "0011"; d4 <= "0001"; -- 1315
    when "0000010100100100" => d1 <= "0110"; d2 <= "0001"; d3 <= "0011"; d4 <= "0001"; -- 1316
    when "0000010100100101" => d1 <= "0111"; d2 <= "0001"; d3 <= "0011"; d4 <= "0001"; -- 1317
    when "0000010100100110" => d1 <= "1000"; d2 <= "0001"; d3 <= "0011"; d4 <= "0001"; -- 1318
    when "0000010100100111" => d1 <= "1001"; d2 <= "0001"; d3 <= "0011"; d4 <= "0001"; -- 1319
    when "0000010100101000" => d1 <= "0000"; d2 <= "0010"; d3 <= "0011"; d4 <= "0001"; -- 1320
    when "0000010100101001" => d1 <= "0001"; d2 <= "0010"; d3 <= "0011"; d4 <= "0001"; -- 1321
    when "0000010100101010" => d1 <= "0010"; d2 <= "0010"; d3 <= "0011"; d4 <= "0001"; -- 1322
    when "0000010100101011" => d1 <= "0011"; d2 <= "0010"; d3 <= "0011"; d4 <= "0001"; -- 1323
    when "0000010100101100" => d1 <= "0100"; d2 <= "0010"; d3 <= "0011"; d4 <= "0001"; -- 1324
    when "0000010100101101" => d1 <= "0101"; d2 <= "0010"; d3 <= "0011"; d4 <= "0001"; -- 1325
    when "0000010100101110" => d1 <= "0110"; d2 <= "0010"; d3 <= "0011"; d4 <= "0001"; -- 1326
    when "0000010100101111" => d1 <= "0111"; d2 <= "0010"; d3 <= "0011"; d4 <= "0001"; -- 1327
    when "0000010100110000" => d1 <= "1000"; d2 <= "0010"; d3 <= "0011"; d4 <= "0001"; -- 1328
    when "0000010100110001" => d1 <= "1001"; d2 <= "0010"; d3 <= "0011"; d4 <= "0001"; -- 1329
    when "0000010100110010" => d1 <= "0000"; d2 <= "0011"; d3 <= "0011"; d4 <= "0001"; -- 1330
    when "0000010100110011" => d1 <= "0001"; d2 <= "0011"; d3 <= "0011"; d4 <= "0001"; -- 1331
    when "0000010100110100" => d1 <= "0010"; d2 <= "0011"; d3 <= "0011"; d4 <= "0001"; -- 1332
    when "0000010100110101" => d1 <= "0011"; d2 <= "0011"; d3 <= "0011"; d4 <= "0001"; -- 1333
    when "0000010100110110" => d1 <= "0100"; d2 <= "0011"; d3 <= "0011"; d4 <= "0001"; -- 1334
    when "0000010100110111" => d1 <= "0101"; d2 <= "0011"; d3 <= "0011"; d4 <= "0001"; -- 1335
    when "0000010100111000" => d1 <= "0110"; d2 <= "0011"; d3 <= "0011"; d4 <= "0001"; -- 1336
    when "0000010100111001" => d1 <= "0111"; d2 <= "0011"; d3 <= "0011"; d4 <= "0001"; -- 1337
    when "0000010100111010" => d1 <= "1000"; d2 <= "0011"; d3 <= "0011"; d4 <= "0001"; -- 1338
    when "0000010100111011" => d1 <= "1001"; d2 <= "0011"; d3 <= "0011"; d4 <= "0001"; -- 1339
    when "0000010100111100" => d1 <= "0000"; d2 <= "0100"; d3 <= "0011"; d4 <= "0001"; -- 1340
    when "0000010100111101" => d1 <= "0001"; d2 <= "0100"; d3 <= "0011"; d4 <= "0001"; -- 1341
    when "0000010100111110" => d1 <= "0010"; d2 <= "0100"; d3 <= "0011"; d4 <= "0001"; -- 1342
    when "0000010100111111" => d1 <= "0011"; d2 <= "0100"; d3 <= "0011"; d4 <= "0001"; -- 1343
    when "0000010101000000" => d1 <= "0100"; d2 <= "0100"; d3 <= "0011"; d4 <= "0001"; -- 1344
    when "0000010101000001" => d1 <= "0101"; d2 <= "0100"; d3 <= "0011"; d4 <= "0001"; -- 1345
    when "0000010101000010" => d1 <= "0110"; d2 <= "0100"; d3 <= "0011"; d4 <= "0001"; -- 1346
    when "0000010101000011" => d1 <= "0111"; d2 <= "0100"; d3 <= "0011"; d4 <= "0001"; -- 1347
    when "0000010101000100" => d1 <= "1000"; d2 <= "0100"; d3 <= "0011"; d4 <= "0001"; -- 1348
    when "0000010101000101" => d1 <= "1001"; d2 <= "0100"; d3 <= "0011"; d4 <= "0001"; -- 1349
    when "0000010101000110" => d1 <= "0000"; d2 <= "0101"; d3 <= "0011"; d4 <= "0001"; -- 1350
    when "0000010101000111" => d1 <= "0001"; d2 <= "0101"; d3 <= "0011"; d4 <= "0001"; -- 1351
    when "0000010101001000" => d1 <= "0010"; d2 <= "0101"; d3 <= "0011"; d4 <= "0001"; -- 1352
    when "0000010101001001" => d1 <= "0011"; d2 <= "0101"; d3 <= "0011"; d4 <= "0001"; -- 1353
    when "0000010101001010" => d1 <= "0100"; d2 <= "0101"; d3 <= "0011"; d4 <= "0001"; -- 1354
    when "0000010101001011" => d1 <= "0101"; d2 <= "0101"; d3 <= "0011"; d4 <= "0001"; -- 1355
    when "0000010101001100" => d1 <= "0110"; d2 <= "0101"; d3 <= "0011"; d4 <= "0001"; -- 1356
    when "0000010101001101" => d1 <= "0111"; d2 <= "0101"; d3 <= "0011"; d4 <= "0001"; -- 1357
    when "0000010101001110" => d1 <= "1000"; d2 <= "0101"; d3 <= "0011"; d4 <= "0001"; -- 1358
    when "0000010101001111" => d1 <= "1001"; d2 <= "0101"; d3 <= "0011"; d4 <= "0001"; -- 1359
    when "0000010101010000" => d1 <= "0000"; d2 <= "0110"; d3 <= "0011"; d4 <= "0001"; -- 1360
    when "0000010101010001" => d1 <= "0001"; d2 <= "0110"; d3 <= "0011"; d4 <= "0001"; -- 1361
    when "0000010101010010" => d1 <= "0010"; d2 <= "0110"; d3 <= "0011"; d4 <= "0001"; -- 1362
    when "0000010101010011" => d1 <= "0011"; d2 <= "0110"; d3 <= "0011"; d4 <= "0001"; -- 1363
    when "0000010101010100" => d1 <= "0100"; d2 <= "0110"; d3 <= "0011"; d4 <= "0001"; -- 1364
    when "0000010101010101" => d1 <= "0101"; d2 <= "0110"; d3 <= "0011"; d4 <= "0001"; -- 1365
    when "0000010101010110" => d1 <= "0110"; d2 <= "0110"; d3 <= "0011"; d4 <= "0001"; -- 1366
    when "0000010101010111" => d1 <= "0111"; d2 <= "0110"; d3 <= "0011"; d4 <= "0001"; -- 1367
    when "0000010101011000" => d1 <= "1000"; d2 <= "0110"; d3 <= "0011"; d4 <= "0001"; -- 1368
    when "0000010101011001" => d1 <= "1001"; d2 <= "0110"; d3 <= "0011"; d4 <= "0001"; -- 1369
    when "0000010101011010" => d1 <= "0000"; d2 <= "0111"; d3 <= "0011"; d4 <= "0001"; -- 1370
    when "0000010101011011" => d1 <= "0001"; d2 <= "0111"; d3 <= "0011"; d4 <= "0001"; -- 1371
    when "0000010101011100" => d1 <= "0010"; d2 <= "0111"; d3 <= "0011"; d4 <= "0001"; -- 1372
    when "0000010101011101" => d1 <= "0011"; d2 <= "0111"; d3 <= "0011"; d4 <= "0001"; -- 1373
    when "0000010101011110" => d1 <= "0100"; d2 <= "0111"; d3 <= "0011"; d4 <= "0001"; -- 1374
    when "0000010101011111" => d1 <= "0101"; d2 <= "0111"; d3 <= "0011"; d4 <= "0001"; -- 1375
    when "0000010101100000" => d1 <= "0110"; d2 <= "0111"; d3 <= "0011"; d4 <= "0001"; -- 1376
    when "0000010101100001" => d1 <= "0111"; d2 <= "0111"; d3 <= "0011"; d4 <= "0001"; -- 1377
    when "0000010101100010" => d1 <= "1000"; d2 <= "0111"; d3 <= "0011"; d4 <= "0001"; -- 1378
    when "0000010101100011" => d1 <= "1001"; d2 <= "0111"; d3 <= "0011"; d4 <= "0001"; -- 1379
    when "0000010101100100" => d1 <= "0000"; d2 <= "1000"; d3 <= "0011"; d4 <= "0001"; -- 1380
    when "0000010101100101" => d1 <= "0001"; d2 <= "1000"; d3 <= "0011"; d4 <= "0001"; -- 1381
    when "0000010101100110" => d1 <= "0010"; d2 <= "1000"; d3 <= "0011"; d4 <= "0001"; -- 1382
    when "0000010101100111" => d1 <= "0011"; d2 <= "1000"; d3 <= "0011"; d4 <= "0001"; -- 1383
    when "0000010101101000" => d1 <= "0100"; d2 <= "1000"; d3 <= "0011"; d4 <= "0001"; -- 1384
    when "0000010101101001" => d1 <= "0101"; d2 <= "1000"; d3 <= "0011"; d4 <= "0001"; -- 1385
    when "0000010101101010" => d1 <= "0110"; d2 <= "1000"; d3 <= "0011"; d4 <= "0001"; -- 1386
    when "0000010101101011" => d1 <= "0111"; d2 <= "1000"; d3 <= "0011"; d4 <= "0001"; -- 1387
    when "0000010101101100" => d1 <= "1000"; d2 <= "1000"; d3 <= "0011"; d4 <= "0001"; -- 1388
    when "0000010101101101" => d1 <= "1001"; d2 <= "1000"; d3 <= "0011"; d4 <= "0001"; -- 1389
    when "0000010101101110" => d1 <= "0000"; d2 <= "1001"; d3 <= "0011"; d4 <= "0001"; -- 1390
    when "0000010101101111" => d1 <= "0001"; d2 <= "1001"; d3 <= "0011"; d4 <= "0001"; -- 1391
    when "0000010101110000" => d1 <= "0010"; d2 <= "1001"; d3 <= "0011"; d4 <= "0001"; -- 1392
    when "0000010101110001" => d1 <= "0011"; d2 <= "1001"; d3 <= "0011"; d4 <= "0001"; -- 1393
    when "0000010101110010" => d1 <= "0100"; d2 <= "1001"; d3 <= "0011"; d4 <= "0001"; -- 1394
    when "0000010101110011" => d1 <= "0101"; d2 <= "1001"; d3 <= "0011"; d4 <= "0001"; -- 1395
    when "0000010101110100" => d1 <= "0110"; d2 <= "1001"; d3 <= "0011"; d4 <= "0001"; -- 1396
    when "0000010101110101" => d1 <= "0111"; d2 <= "1001"; d3 <= "0011"; d4 <= "0001"; -- 1397
    when "0000010101110110" => d1 <= "1000"; d2 <= "1001"; d3 <= "0011"; d4 <= "0001"; -- 1398
    when "0000010101110111" => d1 <= "1001"; d2 <= "1001"; d3 <= "0011"; d4 <= "0001"; -- 1399
    when "0000010101111000" => d1 <= "0000"; d2 <= "0000"; d3 <= "0100"; d4 <= "0001"; -- 1400
    when "0000010101111001" => d1 <= "0001"; d2 <= "0000"; d3 <= "0100"; d4 <= "0001"; -- 1401
    when "0000010101111010" => d1 <= "0010"; d2 <= "0000"; d3 <= "0100"; d4 <= "0001"; -- 1402
    when "0000010101111011" => d1 <= "0011"; d2 <= "0000"; d3 <= "0100"; d4 <= "0001"; -- 1403
    when "0000010101111100" => d1 <= "0100"; d2 <= "0000"; d3 <= "0100"; d4 <= "0001"; -- 1404
    when "0000010101111101" => d1 <= "0101"; d2 <= "0000"; d3 <= "0100"; d4 <= "0001"; -- 1405
    when "0000010101111110" => d1 <= "0110"; d2 <= "0000"; d3 <= "0100"; d4 <= "0001"; -- 1406
    when "0000010101111111" => d1 <= "0111"; d2 <= "0000"; d3 <= "0100"; d4 <= "0001"; -- 1407
    when "0000010110000000" => d1 <= "1000"; d2 <= "0000"; d3 <= "0100"; d4 <= "0001"; -- 1408
    when "0000010110000001" => d1 <= "1001"; d2 <= "0000"; d3 <= "0100"; d4 <= "0001"; -- 1409
    when "0000010110000010" => d1 <= "0000"; d2 <= "0001"; d3 <= "0100"; d4 <= "0001"; -- 1410
    when "0000010110000011" => d1 <= "0001"; d2 <= "0001"; d3 <= "0100"; d4 <= "0001"; -- 1411
    when "0000010110000100" => d1 <= "0010"; d2 <= "0001"; d3 <= "0100"; d4 <= "0001"; -- 1412
    when "0000010110000101" => d1 <= "0011"; d2 <= "0001"; d3 <= "0100"; d4 <= "0001"; -- 1413
    when "0000010110000110" => d1 <= "0100"; d2 <= "0001"; d3 <= "0100"; d4 <= "0001"; -- 1414
    when "0000010110000111" => d1 <= "0101"; d2 <= "0001"; d3 <= "0100"; d4 <= "0001"; -- 1415
    when "0000010110001000" => d1 <= "0110"; d2 <= "0001"; d3 <= "0100"; d4 <= "0001"; -- 1416
    when "0000010110001001" => d1 <= "0111"; d2 <= "0001"; d3 <= "0100"; d4 <= "0001"; -- 1417
    when "0000010110001010" => d1 <= "1000"; d2 <= "0001"; d3 <= "0100"; d4 <= "0001"; -- 1418
    when "0000010110001011" => d1 <= "1001"; d2 <= "0001"; d3 <= "0100"; d4 <= "0001"; -- 1419
    when "0000010110001100" => d1 <= "0000"; d2 <= "0010"; d3 <= "0100"; d4 <= "0001"; -- 1420
    when "0000010110001101" => d1 <= "0001"; d2 <= "0010"; d3 <= "0100"; d4 <= "0001"; -- 1421
    when "0000010110001110" => d1 <= "0010"; d2 <= "0010"; d3 <= "0100"; d4 <= "0001"; -- 1422
    when "0000010110001111" => d1 <= "0011"; d2 <= "0010"; d3 <= "0100"; d4 <= "0001"; -- 1423
    when "0000010110010000" => d1 <= "0100"; d2 <= "0010"; d3 <= "0100"; d4 <= "0001"; -- 1424
    when "0000010110010001" => d1 <= "0101"; d2 <= "0010"; d3 <= "0100"; d4 <= "0001"; -- 1425
    when "0000010110010010" => d1 <= "0110"; d2 <= "0010"; d3 <= "0100"; d4 <= "0001"; -- 1426
    when "0000010110010011" => d1 <= "0111"; d2 <= "0010"; d3 <= "0100"; d4 <= "0001"; -- 1427
    when "0000010110010100" => d1 <= "1000"; d2 <= "0010"; d3 <= "0100"; d4 <= "0001"; -- 1428
    when "0000010110010101" => d1 <= "1001"; d2 <= "0010"; d3 <= "0100"; d4 <= "0001"; -- 1429
    when "0000010110010110" => d1 <= "0000"; d2 <= "0011"; d3 <= "0100"; d4 <= "0001"; -- 1430
    when "0000010110010111" => d1 <= "0001"; d2 <= "0011"; d3 <= "0100"; d4 <= "0001"; -- 1431
    when "0000010110011000" => d1 <= "0010"; d2 <= "0011"; d3 <= "0100"; d4 <= "0001"; -- 1432
    when "0000010110011001" => d1 <= "0011"; d2 <= "0011"; d3 <= "0100"; d4 <= "0001"; -- 1433
    when "0000010110011010" => d1 <= "0100"; d2 <= "0011"; d3 <= "0100"; d4 <= "0001"; -- 1434
    when "0000010110011011" => d1 <= "0101"; d2 <= "0011"; d3 <= "0100"; d4 <= "0001"; -- 1435
    when "0000010110011100" => d1 <= "0110"; d2 <= "0011"; d3 <= "0100"; d4 <= "0001"; -- 1436
    when "0000010110011101" => d1 <= "0111"; d2 <= "0011"; d3 <= "0100"; d4 <= "0001"; -- 1437
    when "0000010110011110" => d1 <= "1000"; d2 <= "0011"; d3 <= "0100"; d4 <= "0001"; -- 1438
    when "0000010110011111" => d1 <= "1001"; d2 <= "0011"; d3 <= "0100"; d4 <= "0001"; -- 1439
    when "0000010110100000" => d1 <= "0000"; d2 <= "0100"; d3 <= "0100"; d4 <= "0001"; -- 1440
    when "0000010110100001" => d1 <= "0001"; d2 <= "0100"; d3 <= "0100"; d4 <= "0001"; -- 1441
    when "0000010110100010" => d1 <= "0010"; d2 <= "0100"; d3 <= "0100"; d4 <= "0001"; -- 1442
    when "0000010110100011" => d1 <= "0011"; d2 <= "0100"; d3 <= "0100"; d4 <= "0001"; -- 1443
    when "0000010110100100" => d1 <= "0100"; d2 <= "0100"; d3 <= "0100"; d4 <= "0001"; -- 1444
    when "0000010110100101" => d1 <= "0101"; d2 <= "0100"; d3 <= "0100"; d4 <= "0001"; -- 1445
    when "0000010110100110" => d1 <= "0110"; d2 <= "0100"; d3 <= "0100"; d4 <= "0001"; -- 1446
    when "0000010110100111" => d1 <= "0111"; d2 <= "0100"; d3 <= "0100"; d4 <= "0001"; -- 1447
    when "0000010110101000" => d1 <= "1000"; d2 <= "0100"; d3 <= "0100"; d4 <= "0001"; -- 1448
    when "0000010110101001" => d1 <= "1001"; d2 <= "0100"; d3 <= "0100"; d4 <= "0001"; -- 1449
    when "0000010110101010" => d1 <= "0000"; d2 <= "0101"; d3 <= "0100"; d4 <= "0001"; -- 1450
    when "0000010110101011" => d1 <= "0001"; d2 <= "0101"; d3 <= "0100"; d4 <= "0001"; -- 1451
    when "0000010110101100" => d1 <= "0010"; d2 <= "0101"; d3 <= "0100"; d4 <= "0001"; -- 1452
    when "0000010110101101" => d1 <= "0011"; d2 <= "0101"; d3 <= "0100"; d4 <= "0001"; -- 1453
    when "0000010110101110" => d1 <= "0100"; d2 <= "0101"; d3 <= "0100"; d4 <= "0001"; -- 1454
    when "0000010110101111" => d1 <= "0101"; d2 <= "0101"; d3 <= "0100"; d4 <= "0001"; -- 1455
    when "0000010110110000" => d1 <= "0110"; d2 <= "0101"; d3 <= "0100"; d4 <= "0001"; -- 1456
    when "0000010110110001" => d1 <= "0111"; d2 <= "0101"; d3 <= "0100"; d4 <= "0001"; -- 1457
    when "0000010110110010" => d1 <= "1000"; d2 <= "0101"; d3 <= "0100"; d4 <= "0001"; -- 1458
    when "0000010110110011" => d1 <= "1001"; d2 <= "0101"; d3 <= "0100"; d4 <= "0001"; -- 1459
    when "0000010110110100" => d1 <= "0000"; d2 <= "0110"; d3 <= "0100"; d4 <= "0001"; -- 1460
    when "0000010110110101" => d1 <= "0001"; d2 <= "0110"; d3 <= "0100"; d4 <= "0001"; -- 1461
    when "0000010110110110" => d1 <= "0010"; d2 <= "0110"; d3 <= "0100"; d4 <= "0001"; -- 1462
    when "0000010110110111" => d1 <= "0011"; d2 <= "0110"; d3 <= "0100"; d4 <= "0001"; -- 1463
    when "0000010110111000" => d1 <= "0100"; d2 <= "0110"; d3 <= "0100"; d4 <= "0001"; -- 1464
    when "0000010110111001" => d1 <= "0101"; d2 <= "0110"; d3 <= "0100"; d4 <= "0001"; -- 1465
    when "0000010110111010" => d1 <= "0110"; d2 <= "0110"; d3 <= "0100"; d4 <= "0001"; -- 1466
    when "0000010110111011" => d1 <= "0111"; d2 <= "0110"; d3 <= "0100"; d4 <= "0001"; -- 1467
    when "0000010110111100" => d1 <= "1000"; d2 <= "0110"; d3 <= "0100"; d4 <= "0001"; -- 1468
    when "0000010110111101" => d1 <= "1001"; d2 <= "0110"; d3 <= "0100"; d4 <= "0001"; -- 1469
    when "0000010110111110" => d1 <= "0000"; d2 <= "0111"; d3 <= "0100"; d4 <= "0001"; -- 1470
    when "0000010110111111" => d1 <= "0001"; d2 <= "0111"; d3 <= "0100"; d4 <= "0001"; -- 1471
    when "0000010111000000" => d1 <= "0010"; d2 <= "0111"; d3 <= "0100"; d4 <= "0001"; -- 1472
    when "0000010111000001" => d1 <= "0011"; d2 <= "0111"; d3 <= "0100"; d4 <= "0001"; -- 1473
    when "0000010111000010" => d1 <= "0100"; d2 <= "0111"; d3 <= "0100"; d4 <= "0001"; -- 1474
    when "0000010111000011" => d1 <= "0101"; d2 <= "0111"; d3 <= "0100"; d4 <= "0001"; -- 1475
    when "0000010111000100" => d1 <= "0110"; d2 <= "0111"; d3 <= "0100"; d4 <= "0001"; -- 1476
    when "0000010111000101" => d1 <= "0111"; d2 <= "0111"; d3 <= "0100"; d4 <= "0001"; -- 1477
    when "0000010111000110" => d1 <= "1000"; d2 <= "0111"; d3 <= "0100"; d4 <= "0001"; -- 1478
    when "0000010111000111" => d1 <= "1001"; d2 <= "0111"; d3 <= "0100"; d4 <= "0001"; -- 1479
    when "0000010111001000" => d1 <= "0000"; d2 <= "1000"; d3 <= "0100"; d4 <= "0001"; -- 1480
    when "0000010111001001" => d1 <= "0001"; d2 <= "1000"; d3 <= "0100"; d4 <= "0001"; -- 1481
    when "0000010111001010" => d1 <= "0010"; d2 <= "1000"; d3 <= "0100"; d4 <= "0001"; -- 1482
    when "0000010111001011" => d1 <= "0011"; d2 <= "1000"; d3 <= "0100"; d4 <= "0001"; -- 1483
    when "0000010111001100" => d1 <= "0100"; d2 <= "1000"; d3 <= "0100"; d4 <= "0001"; -- 1484
    when "0000010111001101" => d1 <= "0101"; d2 <= "1000"; d3 <= "0100"; d4 <= "0001"; -- 1485
    when "0000010111001110" => d1 <= "0110"; d2 <= "1000"; d3 <= "0100"; d4 <= "0001"; -- 1486
    when "0000010111001111" => d1 <= "0111"; d2 <= "1000"; d3 <= "0100"; d4 <= "0001"; -- 1487
    when "0000010111010000" => d1 <= "1000"; d2 <= "1000"; d3 <= "0100"; d4 <= "0001"; -- 1488
    when "0000010111010001" => d1 <= "1001"; d2 <= "1000"; d3 <= "0100"; d4 <= "0001"; -- 1489
    when "0000010111010010" => d1 <= "0000"; d2 <= "1001"; d3 <= "0100"; d4 <= "0001"; -- 1490
    when "0000010111010011" => d1 <= "0001"; d2 <= "1001"; d3 <= "0100"; d4 <= "0001"; -- 1491
    when "0000010111010100" => d1 <= "0010"; d2 <= "1001"; d3 <= "0100"; d4 <= "0001"; -- 1492
    when "0000010111010101" => d1 <= "0011"; d2 <= "1001"; d3 <= "0100"; d4 <= "0001"; -- 1493
    when "0000010111010110" => d1 <= "0100"; d2 <= "1001"; d3 <= "0100"; d4 <= "0001"; -- 1494
    when "0000010111010111" => d1 <= "0101"; d2 <= "1001"; d3 <= "0100"; d4 <= "0001"; -- 1495
    when "0000010111011000" => d1 <= "0110"; d2 <= "1001"; d3 <= "0100"; d4 <= "0001"; -- 1496
    when "0000010111011001" => d1 <= "0111"; d2 <= "1001"; d3 <= "0100"; d4 <= "0001"; -- 1497
    when "0000010111011010" => d1 <= "1000"; d2 <= "1001"; d3 <= "0100"; d4 <= "0001"; -- 1498
    when "0000010111011011" => d1 <= "1001"; d2 <= "1001"; d3 <= "0100"; d4 <= "0001"; -- 1499
    when "0000010111011100" => d1 <= "0000"; d2 <= "0000"; d3 <= "0101"; d4 <= "0001"; -- 1500
    when "0000010111011101" => d1 <= "0001"; d2 <= "0000"; d3 <= "0101"; d4 <= "0001"; -- 1501
    when "0000010111011110" => d1 <= "0010"; d2 <= "0000"; d3 <= "0101"; d4 <= "0001"; -- 1502
    when "0000010111011111" => d1 <= "0011"; d2 <= "0000"; d3 <= "0101"; d4 <= "0001"; -- 1503
    when "0000010111100000" => d1 <= "0100"; d2 <= "0000"; d3 <= "0101"; d4 <= "0001"; -- 1504
    when "0000010111100001" => d1 <= "0101"; d2 <= "0000"; d3 <= "0101"; d4 <= "0001"; -- 1505
    when "0000010111100010" => d1 <= "0110"; d2 <= "0000"; d3 <= "0101"; d4 <= "0001"; -- 1506
    when "0000010111100011" => d1 <= "0111"; d2 <= "0000"; d3 <= "0101"; d4 <= "0001"; -- 1507
    when "0000010111100100" => d1 <= "1000"; d2 <= "0000"; d3 <= "0101"; d4 <= "0001"; -- 1508
    when "0000010111100101" => d1 <= "1001"; d2 <= "0000"; d3 <= "0101"; d4 <= "0001"; -- 1509
    when "0000010111100110" => d1 <= "0000"; d2 <= "0001"; d3 <= "0101"; d4 <= "0001"; -- 1510
    when "0000010111100111" => d1 <= "0001"; d2 <= "0001"; d3 <= "0101"; d4 <= "0001"; -- 1511
    when "0000010111101000" => d1 <= "0010"; d2 <= "0001"; d3 <= "0101"; d4 <= "0001"; -- 1512
    when "0000010111101001" => d1 <= "0011"; d2 <= "0001"; d3 <= "0101"; d4 <= "0001"; -- 1513
    when "0000010111101010" => d1 <= "0100"; d2 <= "0001"; d3 <= "0101"; d4 <= "0001"; -- 1514
    when "0000010111101011" => d1 <= "0101"; d2 <= "0001"; d3 <= "0101"; d4 <= "0001"; -- 1515
    when "0000010111101100" => d1 <= "0110"; d2 <= "0001"; d3 <= "0101"; d4 <= "0001"; -- 1516
    when "0000010111101101" => d1 <= "0111"; d2 <= "0001"; d3 <= "0101"; d4 <= "0001"; -- 1517
    when "0000010111101110" => d1 <= "1000"; d2 <= "0001"; d3 <= "0101"; d4 <= "0001"; -- 1518
    when "0000010111101111" => d1 <= "1001"; d2 <= "0001"; d3 <= "0101"; d4 <= "0001"; -- 1519
    when "0000010111110000" => d1 <= "0000"; d2 <= "0010"; d3 <= "0101"; d4 <= "0001"; -- 1520
    when "0000010111110001" => d1 <= "0001"; d2 <= "0010"; d3 <= "0101"; d4 <= "0001"; -- 1521
    when "0000010111110010" => d1 <= "0010"; d2 <= "0010"; d3 <= "0101"; d4 <= "0001"; -- 1522
    when "0000010111110011" => d1 <= "0011"; d2 <= "0010"; d3 <= "0101"; d4 <= "0001"; -- 1523
    when "0000010111110100" => d1 <= "0100"; d2 <= "0010"; d3 <= "0101"; d4 <= "0001"; -- 1524
    when "0000010111110101" => d1 <= "0101"; d2 <= "0010"; d3 <= "0101"; d4 <= "0001"; -- 1525
    when "0000010111110110" => d1 <= "0110"; d2 <= "0010"; d3 <= "0101"; d4 <= "0001"; -- 1526
    when "0000010111110111" => d1 <= "0111"; d2 <= "0010"; d3 <= "0101"; d4 <= "0001"; -- 1527
    when "0000010111111000" => d1 <= "1000"; d2 <= "0010"; d3 <= "0101"; d4 <= "0001"; -- 1528
    when "0000010111111001" => d1 <= "1001"; d2 <= "0010"; d3 <= "0101"; d4 <= "0001"; -- 1529
    when "0000010111111010" => d1 <= "0000"; d2 <= "0011"; d3 <= "0101"; d4 <= "0001"; -- 1530
    when "0000010111111011" => d1 <= "0001"; d2 <= "0011"; d3 <= "0101"; d4 <= "0001"; -- 1531
    when "0000010111111100" => d1 <= "0010"; d2 <= "0011"; d3 <= "0101"; d4 <= "0001"; -- 1532
    when "0000010111111101" => d1 <= "0011"; d2 <= "0011"; d3 <= "0101"; d4 <= "0001"; -- 1533
    when "0000010111111110" => d1 <= "0100"; d2 <= "0011"; d3 <= "0101"; d4 <= "0001"; -- 1534
    when "0000010111111111" => d1 <= "0101"; d2 <= "0011"; d3 <= "0101"; d4 <= "0001"; -- 1535
    when "0000011000000000" => d1 <= "0110"; d2 <= "0011"; d3 <= "0101"; d4 <= "0001"; -- 1536
    when "0000011000000001" => d1 <= "0111"; d2 <= "0011"; d3 <= "0101"; d4 <= "0001"; -- 1537
    when "0000011000000010" => d1 <= "1000"; d2 <= "0011"; d3 <= "0101"; d4 <= "0001"; -- 1538
    when "0000011000000011" => d1 <= "1001"; d2 <= "0011"; d3 <= "0101"; d4 <= "0001"; -- 1539
    when "0000011000000100" => d1 <= "0000"; d2 <= "0100"; d3 <= "0101"; d4 <= "0001"; -- 1540
    when "0000011000000101" => d1 <= "0001"; d2 <= "0100"; d3 <= "0101"; d4 <= "0001"; -- 1541
    when "0000011000000110" => d1 <= "0010"; d2 <= "0100"; d3 <= "0101"; d4 <= "0001"; -- 1542
    when "0000011000000111" => d1 <= "0011"; d2 <= "0100"; d3 <= "0101"; d4 <= "0001"; -- 1543
    when "0000011000001000" => d1 <= "0100"; d2 <= "0100"; d3 <= "0101"; d4 <= "0001"; -- 1544
    when "0000011000001001" => d1 <= "0101"; d2 <= "0100"; d3 <= "0101"; d4 <= "0001"; -- 1545
    when "0000011000001010" => d1 <= "0110"; d2 <= "0100"; d3 <= "0101"; d4 <= "0001"; -- 1546
    when "0000011000001011" => d1 <= "0111"; d2 <= "0100"; d3 <= "0101"; d4 <= "0001"; -- 1547
    when "0000011000001100" => d1 <= "1000"; d2 <= "0100"; d3 <= "0101"; d4 <= "0001"; -- 1548
    when "0000011000001101" => d1 <= "1001"; d2 <= "0100"; d3 <= "0101"; d4 <= "0001"; -- 1549
    when "0000011000001110" => d1 <= "0000"; d2 <= "0101"; d3 <= "0101"; d4 <= "0001"; -- 1550
    when "0000011000001111" => d1 <= "0001"; d2 <= "0101"; d3 <= "0101"; d4 <= "0001"; -- 1551
    when "0000011000010000" => d1 <= "0010"; d2 <= "0101"; d3 <= "0101"; d4 <= "0001"; -- 1552
    when "0000011000010001" => d1 <= "0011"; d2 <= "0101"; d3 <= "0101"; d4 <= "0001"; -- 1553
    when "0000011000010010" => d1 <= "0100"; d2 <= "0101"; d3 <= "0101"; d4 <= "0001"; -- 1554
    when "0000011000010011" => d1 <= "0101"; d2 <= "0101"; d3 <= "0101"; d4 <= "0001"; -- 1555
    when "0000011000010100" => d1 <= "0110"; d2 <= "0101"; d3 <= "0101"; d4 <= "0001"; -- 1556
    when "0000011000010101" => d1 <= "0111"; d2 <= "0101"; d3 <= "0101"; d4 <= "0001"; -- 1557
    when "0000011000010110" => d1 <= "1000"; d2 <= "0101"; d3 <= "0101"; d4 <= "0001"; -- 1558
    when "0000011000010111" => d1 <= "1001"; d2 <= "0101"; d3 <= "0101"; d4 <= "0001"; -- 1559
    when "0000011000011000" => d1 <= "0000"; d2 <= "0110"; d3 <= "0101"; d4 <= "0001"; -- 1560
    when "0000011000011001" => d1 <= "0001"; d2 <= "0110"; d3 <= "0101"; d4 <= "0001"; -- 1561
    when "0000011000011010" => d1 <= "0010"; d2 <= "0110"; d3 <= "0101"; d4 <= "0001"; -- 1562
    when "0000011000011011" => d1 <= "0011"; d2 <= "0110"; d3 <= "0101"; d4 <= "0001"; -- 1563
    when "0000011000011100" => d1 <= "0100"; d2 <= "0110"; d3 <= "0101"; d4 <= "0001"; -- 1564
    when "0000011000011101" => d1 <= "0101"; d2 <= "0110"; d3 <= "0101"; d4 <= "0001"; -- 1565
    when "0000011000011110" => d1 <= "0110"; d2 <= "0110"; d3 <= "0101"; d4 <= "0001"; -- 1566
    when "0000011000011111" => d1 <= "0111"; d2 <= "0110"; d3 <= "0101"; d4 <= "0001"; -- 1567
    when "0000011000100000" => d1 <= "1000"; d2 <= "0110"; d3 <= "0101"; d4 <= "0001"; -- 1568
    when "0000011000100001" => d1 <= "1001"; d2 <= "0110"; d3 <= "0101"; d4 <= "0001"; -- 1569
    when "0000011000100010" => d1 <= "0000"; d2 <= "0111"; d3 <= "0101"; d4 <= "0001"; -- 1570
    when "0000011000100011" => d1 <= "0001"; d2 <= "0111"; d3 <= "0101"; d4 <= "0001"; -- 1571
    when "0000011000100100" => d1 <= "0010"; d2 <= "0111"; d3 <= "0101"; d4 <= "0001"; -- 1572
    when "0000011000100101" => d1 <= "0011"; d2 <= "0111"; d3 <= "0101"; d4 <= "0001"; -- 1573
    when "0000011000100110" => d1 <= "0100"; d2 <= "0111"; d3 <= "0101"; d4 <= "0001"; -- 1574
    when "0000011000100111" => d1 <= "0101"; d2 <= "0111"; d3 <= "0101"; d4 <= "0001"; -- 1575
    when "0000011000101000" => d1 <= "0110"; d2 <= "0111"; d3 <= "0101"; d4 <= "0001"; -- 1576
    when "0000011000101001" => d1 <= "0111"; d2 <= "0111"; d3 <= "0101"; d4 <= "0001"; -- 1577
    when "0000011000101010" => d1 <= "1000"; d2 <= "0111"; d3 <= "0101"; d4 <= "0001"; -- 1578
    when "0000011000101011" => d1 <= "1001"; d2 <= "0111"; d3 <= "0101"; d4 <= "0001"; -- 1579
    when "0000011000101100" => d1 <= "0000"; d2 <= "1000"; d3 <= "0101"; d4 <= "0001"; -- 1580
    when "0000011000101101" => d1 <= "0001"; d2 <= "1000"; d3 <= "0101"; d4 <= "0001"; -- 1581
    when "0000011000101110" => d1 <= "0010"; d2 <= "1000"; d3 <= "0101"; d4 <= "0001"; -- 1582
    when "0000011000101111" => d1 <= "0011"; d2 <= "1000"; d3 <= "0101"; d4 <= "0001"; -- 1583
    when "0000011000110000" => d1 <= "0100"; d2 <= "1000"; d3 <= "0101"; d4 <= "0001"; -- 1584
    when "0000011000110001" => d1 <= "0101"; d2 <= "1000"; d3 <= "0101"; d4 <= "0001"; -- 1585
    when "0000011000110010" => d1 <= "0110"; d2 <= "1000"; d3 <= "0101"; d4 <= "0001"; -- 1586
    when "0000011000110011" => d1 <= "0111"; d2 <= "1000"; d3 <= "0101"; d4 <= "0001"; -- 1587
    when "0000011000110100" => d1 <= "1000"; d2 <= "1000"; d3 <= "0101"; d4 <= "0001"; -- 1588
    when "0000011000110101" => d1 <= "1001"; d2 <= "1000"; d3 <= "0101"; d4 <= "0001"; -- 1589
    when "0000011000110110" => d1 <= "0000"; d2 <= "1001"; d3 <= "0101"; d4 <= "0001"; -- 1590
    when "0000011000110111" => d1 <= "0001"; d2 <= "1001"; d3 <= "0101"; d4 <= "0001"; -- 1591
    when "0000011000111000" => d1 <= "0010"; d2 <= "1001"; d3 <= "0101"; d4 <= "0001"; -- 1592
    when "0000011000111001" => d1 <= "0011"; d2 <= "1001"; d3 <= "0101"; d4 <= "0001"; -- 1593
    when "0000011000111010" => d1 <= "0100"; d2 <= "1001"; d3 <= "0101"; d4 <= "0001"; -- 1594
    when "0000011000111011" => d1 <= "0101"; d2 <= "1001"; d3 <= "0101"; d4 <= "0001"; -- 1595
    when "0000011000111100" => d1 <= "0110"; d2 <= "1001"; d3 <= "0101"; d4 <= "0001"; -- 1596
    when "0000011000111101" => d1 <= "0111"; d2 <= "1001"; d3 <= "0101"; d4 <= "0001"; -- 1597
    when "0000011000111110" => d1 <= "1000"; d2 <= "1001"; d3 <= "0101"; d4 <= "0001"; -- 1598
    when "0000011000111111" => d1 <= "1001"; d2 <= "1001"; d3 <= "0101"; d4 <= "0001"; -- 1599
    when "0000011001000000" => d1 <= "0000"; d2 <= "0000"; d3 <= "0110"; d4 <= "0001"; -- 1600
    when "0000011001000001" => d1 <= "0001"; d2 <= "0000"; d3 <= "0110"; d4 <= "0001"; -- 1601
    when "0000011001000010" => d1 <= "0010"; d2 <= "0000"; d3 <= "0110"; d4 <= "0001"; -- 1602
    when "0000011001000011" => d1 <= "0011"; d2 <= "0000"; d3 <= "0110"; d4 <= "0001"; -- 1603
    when "0000011001000100" => d1 <= "0100"; d2 <= "0000"; d3 <= "0110"; d4 <= "0001"; -- 1604
    when "0000011001000101" => d1 <= "0101"; d2 <= "0000"; d3 <= "0110"; d4 <= "0001"; -- 1605
    when "0000011001000110" => d1 <= "0110"; d2 <= "0000"; d3 <= "0110"; d4 <= "0001"; -- 1606
    when "0000011001000111" => d1 <= "0111"; d2 <= "0000"; d3 <= "0110"; d4 <= "0001"; -- 1607
    when "0000011001001000" => d1 <= "1000"; d2 <= "0000"; d3 <= "0110"; d4 <= "0001"; -- 1608
    when "0000011001001001" => d1 <= "1001"; d2 <= "0000"; d3 <= "0110"; d4 <= "0001"; -- 1609
    when "0000011001001010" => d1 <= "0000"; d2 <= "0001"; d3 <= "0110"; d4 <= "0001"; -- 1610
    when "0000011001001011" => d1 <= "0001"; d2 <= "0001"; d3 <= "0110"; d4 <= "0001"; -- 1611
    when "0000011001001100" => d1 <= "0010"; d2 <= "0001"; d3 <= "0110"; d4 <= "0001"; -- 1612
    when "0000011001001101" => d1 <= "0011"; d2 <= "0001"; d3 <= "0110"; d4 <= "0001"; -- 1613
    when "0000011001001110" => d1 <= "0100"; d2 <= "0001"; d3 <= "0110"; d4 <= "0001"; -- 1614
    when "0000011001001111" => d1 <= "0101"; d2 <= "0001"; d3 <= "0110"; d4 <= "0001"; -- 1615
    when "0000011001010000" => d1 <= "0110"; d2 <= "0001"; d3 <= "0110"; d4 <= "0001"; -- 1616
    when "0000011001010001" => d1 <= "0111"; d2 <= "0001"; d3 <= "0110"; d4 <= "0001"; -- 1617
    when "0000011001010010" => d1 <= "1000"; d2 <= "0001"; d3 <= "0110"; d4 <= "0001"; -- 1618
    when "0000011001010011" => d1 <= "1001"; d2 <= "0001"; d3 <= "0110"; d4 <= "0001"; -- 1619
    when "0000011001010100" => d1 <= "0000"; d2 <= "0010"; d3 <= "0110"; d4 <= "0001"; -- 1620
    when "0000011001010101" => d1 <= "0001"; d2 <= "0010"; d3 <= "0110"; d4 <= "0001"; -- 1621
    when "0000011001010110" => d1 <= "0010"; d2 <= "0010"; d3 <= "0110"; d4 <= "0001"; -- 1622
    when "0000011001010111" => d1 <= "0011"; d2 <= "0010"; d3 <= "0110"; d4 <= "0001"; -- 1623
    when "0000011001011000" => d1 <= "0100"; d2 <= "0010"; d3 <= "0110"; d4 <= "0001"; -- 1624
    when "0000011001011001" => d1 <= "0101"; d2 <= "0010"; d3 <= "0110"; d4 <= "0001"; -- 1625
    when "0000011001011010" => d1 <= "0110"; d2 <= "0010"; d3 <= "0110"; d4 <= "0001"; -- 1626
    when "0000011001011011" => d1 <= "0111"; d2 <= "0010"; d3 <= "0110"; d4 <= "0001"; -- 1627
    when "0000011001011100" => d1 <= "1000"; d2 <= "0010"; d3 <= "0110"; d4 <= "0001"; -- 1628
    when "0000011001011101" => d1 <= "1001"; d2 <= "0010"; d3 <= "0110"; d4 <= "0001"; -- 1629
    when "0000011001011110" => d1 <= "0000"; d2 <= "0011"; d3 <= "0110"; d4 <= "0001"; -- 1630
    when "0000011001011111" => d1 <= "0001"; d2 <= "0011"; d3 <= "0110"; d4 <= "0001"; -- 1631
    when "0000011001100000" => d1 <= "0010"; d2 <= "0011"; d3 <= "0110"; d4 <= "0001"; -- 1632
    when "0000011001100001" => d1 <= "0011"; d2 <= "0011"; d3 <= "0110"; d4 <= "0001"; -- 1633
    when "0000011001100010" => d1 <= "0100"; d2 <= "0011"; d3 <= "0110"; d4 <= "0001"; -- 1634
    when "0000011001100011" => d1 <= "0101"; d2 <= "0011"; d3 <= "0110"; d4 <= "0001"; -- 1635
    when "0000011001100100" => d1 <= "0110"; d2 <= "0011"; d3 <= "0110"; d4 <= "0001"; -- 1636
    when "0000011001100101" => d1 <= "0111"; d2 <= "0011"; d3 <= "0110"; d4 <= "0001"; -- 1637
    when "0000011001100110" => d1 <= "1000"; d2 <= "0011"; d3 <= "0110"; d4 <= "0001"; -- 1638
    when "0000011001100111" => d1 <= "1001"; d2 <= "0011"; d3 <= "0110"; d4 <= "0001"; -- 1639
    when "0000011001101000" => d1 <= "0000"; d2 <= "0100"; d3 <= "0110"; d4 <= "0001"; -- 1640
    when "0000011001101001" => d1 <= "0001"; d2 <= "0100"; d3 <= "0110"; d4 <= "0001"; -- 1641
    when "0000011001101010" => d1 <= "0010"; d2 <= "0100"; d3 <= "0110"; d4 <= "0001"; -- 1642
    when "0000011001101011" => d1 <= "0011"; d2 <= "0100"; d3 <= "0110"; d4 <= "0001"; -- 1643
    when "0000011001101100" => d1 <= "0100"; d2 <= "0100"; d3 <= "0110"; d4 <= "0001"; -- 1644
    when "0000011001101101" => d1 <= "0101"; d2 <= "0100"; d3 <= "0110"; d4 <= "0001"; -- 1645
    when "0000011001101110" => d1 <= "0110"; d2 <= "0100"; d3 <= "0110"; d4 <= "0001"; -- 1646
    when "0000011001101111" => d1 <= "0111"; d2 <= "0100"; d3 <= "0110"; d4 <= "0001"; -- 1647
    when "0000011001110000" => d1 <= "1000"; d2 <= "0100"; d3 <= "0110"; d4 <= "0001"; -- 1648
    when "0000011001110001" => d1 <= "1001"; d2 <= "0100"; d3 <= "0110"; d4 <= "0001"; -- 1649
    when "0000011001110010" => d1 <= "0000"; d2 <= "0101"; d3 <= "0110"; d4 <= "0001"; -- 1650
    when "0000011001110011" => d1 <= "0001"; d2 <= "0101"; d3 <= "0110"; d4 <= "0001"; -- 1651
    when "0000011001110100" => d1 <= "0010"; d2 <= "0101"; d3 <= "0110"; d4 <= "0001"; -- 1652
    when "0000011001110101" => d1 <= "0011"; d2 <= "0101"; d3 <= "0110"; d4 <= "0001"; -- 1653
    when "0000011001110110" => d1 <= "0100"; d2 <= "0101"; d3 <= "0110"; d4 <= "0001"; -- 1654
    when "0000011001110111" => d1 <= "0101"; d2 <= "0101"; d3 <= "0110"; d4 <= "0001"; -- 1655
    when "0000011001111000" => d1 <= "0110"; d2 <= "0101"; d3 <= "0110"; d4 <= "0001"; -- 1656
    when "0000011001111001" => d1 <= "0111"; d2 <= "0101"; d3 <= "0110"; d4 <= "0001"; -- 1657
    when "0000011001111010" => d1 <= "1000"; d2 <= "0101"; d3 <= "0110"; d4 <= "0001"; -- 1658
    when "0000011001111011" => d1 <= "1001"; d2 <= "0101"; d3 <= "0110"; d4 <= "0001"; -- 1659
    when "0000011001111100" => d1 <= "0000"; d2 <= "0110"; d3 <= "0110"; d4 <= "0001"; -- 1660
    when "0000011001111101" => d1 <= "0001"; d2 <= "0110"; d3 <= "0110"; d4 <= "0001"; -- 1661
    when "0000011001111110" => d1 <= "0010"; d2 <= "0110"; d3 <= "0110"; d4 <= "0001"; -- 1662
    when "0000011001111111" => d1 <= "0011"; d2 <= "0110"; d3 <= "0110"; d4 <= "0001"; -- 1663
    when "0000011010000000" => d1 <= "0100"; d2 <= "0110"; d3 <= "0110"; d4 <= "0001"; -- 1664
    when "0000011010000001" => d1 <= "0101"; d2 <= "0110"; d3 <= "0110"; d4 <= "0001"; -- 1665
    when "0000011010000010" => d1 <= "0110"; d2 <= "0110"; d3 <= "0110"; d4 <= "0001"; -- 1666
    when "0000011010000011" => d1 <= "0111"; d2 <= "0110"; d3 <= "0110"; d4 <= "0001"; -- 1667
    when "0000011010000100" => d1 <= "1000"; d2 <= "0110"; d3 <= "0110"; d4 <= "0001"; -- 1668
    when "0000011010000101" => d1 <= "1001"; d2 <= "0110"; d3 <= "0110"; d4 <= "0001"; -- 1669
    when "0000011010000110" => d1 <= "0000"; d2 <= "0111"; d3 <= "0110"; d4 <= "0001"; -- 1670
    when "0000011010000111" => d1 <= "0001"; d2 <= "0111"; d3 <= "0110"; d4 <= "0001"; -- 1671
    when "0000011010001000" => d1 <= "0010"; d2 <= "0111"; d3 <= "0110"; d4 <= "0001"; -- 1672
    when "0000011010001001" => d1 <= "0011"; d2 <= "0111"; d3 <= "0110"; d4 <= "0001"; -- 1673
    when "0000011010001010" => d1 <= "0100"; d2 <= "0111"; d3 <= "0110"; d4 <= "0001"; -- 1674
    when "0000011010001011" => d1 <= "0101"; d2 <= "0111"; d3 <= "0110"; d4 <= "0001"; -- 1675
    when "0000011010001100" => d1 <= "0110"; d2 <= "0111"; d3 <= "0110"; d4 <= "0001"; -- 1676
    when "0000011010001101" => d1 <= "0111"; d2 <= "0111"; d3 <= "0110"; d4 <= "0001"; -- 1677
    when "0000011010001110" => d1 <= "1000"; d2 <= "0111"; d3 <= "0110"; d4 <= "0001"; -- 1678
    when "0000011010001111" => d1 <= "1001"; d2 <= "0111"; d3 <= "0110"; d4 <= "0001"; -- 1679
    when "0000011010010000" => d1 <= "0000"; d2 <= "1000"; d3 <= "0110"; d4 <= "0001"; -- 1680
    when "0000011010010001" => d1 <= "0001"; d2 <= "1000"; d3 <= "0110"; d4 <= "0001"; -- 1681
    when "0000011010010010" => d1 <= "0010"; d2 <= "1000"; d3 <= "0110"; d4 <= "0001"; -- 1682
    when "0000011010010011" => d1 <= "0011"; d2 <= "1000"; d3 <= "0110"; d4 <= "0001"; -- 1683
    when "0000011010010100" => d1 <= "0100"; d2 <= "1000"; d3 <= "0110"; d4 <= "0001"; -- 1684
    when "0000011010010101" => d1 <= "0101"; d2 <= "1000"; d3 <= "0110"; d4 <= "0001"; -- 1685
    when "0000011010010110" => d1 <= "0110"; d2 <= "1000"; d3 <= "0110"; d4 <= "0001"; -- 1686
    when "0000011010010111" => d1 <= "0111"; d2 <= "1000"; d3 <= "0110"; d4 <= "0001"; -- 1687
    when "0000011010011000" => d1 <= "1000"; d2 <= "1000"; d3 <= "0110"; d4 <= "0001"; -- 1688
    when "0000011010011001" => d1 <= "1001"; d2 <= "1000"; d3 <= "0110"; d4 <= "0001"; -- 1689
    when "0000011010011010" => d1 <= "0000"; d2 <= "1001"; d3 <= "0110"; d4 <= "0001"; -- 1690
    when "0000011010011011" => d1 <= "0001"; d2 <= "1001"; d3 <= "0110"; d4 <= "0001"; -- 1691
    when "0000011010011100" => d1 <= "0010"; d2 <= "1001"; d3 <= "0110"; d4 <= "0001"; -- 1692
    when "0000011010011101" => d1 <= "0011"; d2 <= "1001"; d3 <= "0110"; d4 <= "0001"; -- 1693
    when "0000011010011110" => d1 <= "0100"; d2 <= "1001"; d3 <= "0110"; d4 <= "0001"; -- 1694
    when "0000011010011111" => d1 <= "0101"; d2 <= "1001"; d3 <= "0110"; d4 <= "0001"; -- 1695
    when "0000011010100000" => d1 <= "0110"; d2 <= "1001"; d3 <= "0110"; d4 <= "0001"; -- 1696
    when "0000011010100001" => d1 <= "0111"; d2 <= "1001"; d3 <= "0110"; d4 <= "0001"; -- 1697
    when "0000011010100010" => d1 <= "1000"; d2 <= "1001"; d3 <= "0110"; d4 <= "0001"; -- 1698
    when "0000011010100011" => d1 <= "1001"; d2 <= "1001"; d3 <= "0110"; d4 <= "0001"; -- 1699
    when "0000011010100100" => d1 <= "0000"; d2 <= "0000"; d3 <= "0111"; d4 <= "0001"; -- 1700
    when "0000011010100101" => d1 <= "0001"; d2 <= "0000"; d3 <= "0111"; d4 <= "0001"; -- 1701
    when "0000011010100110" => d1 <= "0010"; d2 <= "0000"; d3 <= "0111"; d4 <= "0001"; -- 1702
    when "0000011010100111" => d1 <= "0011"; d2 <= "0000"; d3 <= "0111"; d4 <= "0001"; -- 1703
    when "0000011010101000" => d1 <= "0100"; d2 <= "0000"; d3 <= "0111"; d4 <= "0001"; -- 1704
    when "0000011010101001" => d1 <= "0101"; d2 <= "0000"; d3 <= "0111"; d4 <= "0001"; -- 1705
    when "0000011010101010" => d1 <= "0110"; d2 <= "0000"; d3 <= "0111"; d4 <= "0001"; -- 1706
    when "0000011010101011" => d1 <= "0111"; d2 <= "0000"; d3 <= "0111"; d4 <= "0001"; -- 1707
    when "0000011010101100" => d1 <= "1000"; d2 <= "0000"; d3 <= "0111"; d4 <= "0001"; -- 1708
    when "0000011010101101" => d1 <= "1001"; d2 <= "0000"; d3 <= "0111"; d4 <= "0001"; -- 1709
    when "0000011010101110" => d1 <= "0000"; d2 <= "0001"; d3 <= "0111"; d4 <= "0001"; -- 1710
    when "0000011010101111" => d1 <= "0001"; d2 <= "0001"; d3 <= "0111"; d4 <= "0001"; -- 1711
    when "0000011010110000" => d1 <= "0010"; d2 <= "0001"; d3 <= "0111"; d4 <= "0001"; -- 1712
    when "0000011010110001" => d1 <= "0011"; d2 <= "0001"; d3 <= "0111"; d4 <= "0001"; -- 1713
    when "0000011010110010" => d1 <= "0100"; d2 <= "0001"; d3 <= "0111"; d4 <= "0001"; -- 1714
    when "0000011010110011" => d1 <= "0101"; d2 <= "0001"; d3 <= "0111"; d4 <= "0001"; -- 1715
    when "0000011010110100" => d1 <= "0110"; d2 <= "0001"; d3 <= "0111"; d4 <= "0001"; -- 1716
    when "0000011010110101" => d1 <= "0111"; d2 <= "0001"; d3 <= "0111"; d4 <= "0001"; -- 1717
    when "0000011010110110" => d1 <= "1000"; d2 <= "0001"; d3 <= "0111"; d4 <= "0001"; -- 1718
    when "0000011010110111" => d1 <= "1001"; d2 <= "0001"; d3 <= "0111"; d4 <= "0001"; -- 1719
    when "0000011010111000" => d1 <= "0000"; d2 <= "0010"; d3 <= "0111"; d4 <= "0001"; -- 1720
    when "0000011010111001" => d1 <= "0001"; d2 <= "0010"; d3 <= "0111"; d4 <= "0001"; -- 1721
    when "0000011010111010" => d1 <= "0010"; d2 <= "0010"; d3 <= "0111"; d4 <= "0001"; -- 1722
    when "0000011010111011" => d1 <= "0011"; d2 <= "0010"; d3 <= "0111"; d4 <= "0001"; -- 1723
    when "0000011010111100" => d1 <= "0100"; d2 <= "0010"; d3 <= "0111"; d4 <= "0001"; -- 1724
    when "0000011010111101" => d1 <= "0101"; d2 <= "0010"; d3 <= "0111"; d4 <= "0001"; -- 1725
    when "0000011010111110" => d1 <= "0110"; d2 <= "0010"; d3 <= "0111"; d4 <= "0001"; -- 1726
    when "0000011010111111" => d1 <= "0111"; d2 <= "0010"; d3 <= "0111"; d4 <= "0001"; -- 1727
    when "0000011011000000" => d1 <= "1000"; d2 <= "0010"; d3 <= "0111"; d4 <= "0001"; -- 1728
    when "0000011011000001" => d1 <= "1001"; d2 <= "0010"; d3 <= "0111"; d4 <= "0001"; -- 1729
    when "0000011011000010" => d1 <= "0000"; d2 <= "0011"; d3 <= "0111"; d4 <= "0001"; -- 1730
    when "0000011011000011" => d1 <= "0001"; d2 <= "0011"; d3 <= "0111"; d4 <= "0001"; -- 1731
    when "0000011011000100" => d1 <= "0010"; d2 <= "0011"; d3 <= "0111"; d4 <= "0001"; -- 1732
    when "0000011011000101" => d1 <= "0011"; d2 <= "0011"; d3 <= "0111"; d4 <= "0001"; -- 1733
    when "0000011011000110" => d1 <= "0100"; d2 <= "0011"; d3 <= "0111"; d4 <= "0001"; -- 1734
    when "0000011011000111" => d1 <= "0101"; d2 <= "0011"; d3 <= "0111"; d4 <= "0001"; -- 1735
    when "0000011011001000" => d1 <= "0110"; d2 <= "0011"; d3 <= "0111"; d4 <= "0001"; -- 1736
    when "0000011011001001" => d1 <= "0111"; d2 <= "0011"; d3 <= "0111"; d4 <= "0001"; -- 1737
    when "0000011011001010" => d1 <= "1000"; d2 <= "0011"; d3 <= "0111"; d4 <= "0001"; -- 1738
    when "0000011011001011" => d1 <= "1001"; d2 <= "0011"; d3 <= "0111"; d4 <= "0001"; -- 1739
    when "0000011011001100" => d1 <= "0000"; d2 <= "0100"; d3 <= "0111"; d4 <= "0001"; -- 1740
    when "0000011011001101" => d1 <= "0001"; d2 <= "0100"; d3 <= "0111"; d4 <= "0001"; -- 1741
    when "0000011011001110" => d1 <= "0010"; d2 <= "0100"; d3 <= "0111"; d4 <= "0001"; -- 1742
    when "0000011011001111" => d1 <= "0011"; d2 <= "0100"; d3 <= "0111"; d4 <= "0001"; -- 1743
    when "0000011011010000" => d1 <= "0100"; d2 <= "0100"; d3 <= "0111"; d4 <= "0001"; -- 1744
    when "0000011011010001" => d1 <= "0101"; d2 <= "0100"; d3 <= "0111"; d4 <= "0001"; -- 1745
    when "0000011011010010" => d1 <= "0110"; d2 <= "0100"; d3 <= "0111"; d4 <= "0001"; -- 1746
    when "0000011011010011" => d1 <= "0111"; d2 <= "0100"; d3 <= "0111"; d4 <= "0001"; -- 1747
    when "0000011011010100" => d1 <= "1000"; d2 <= "0100"; d3 <= "0111"; d4 <= "0001"; -- 1748
    when "0000011011010101" => d1 <= "1001"; d2 <= "0100"; d3 <= "0111"; d4 <= "0001"; -- 1749
    when "0000011011010110" => d1 <= "0000"; d2 <= "0101"; d3 <= "0111"; d4 <= "0001"; -- 1750
    when "0000011011010111" => d1 <= "0001"; d2 <= "0101"; d3 <= "0111"; d4 <= "0001"; -- 1751
    when "0000011011011000" => d1 <= "0010"; d2 <= "0101"; d3 <= "0111"; d4 <= "0001"; -- 1752
    when "0000011011011001" => d1 <= "0011"; d2 <= "0101"; d3 <= "0111"; d4 <= "0001"; -- 1753
    when "0000011011011010" => d1 <= "0100"; d2 <= "0101"; d3 <= "0111"; d4 <= "0001"; -- 1754
    when "0000011011011011" => d1 <= "0101"; d2 <= "0101"; d3 <= "0111"; d4 <= "0001"; -- 1755
    when "0000011011011100" => d1 <= "0110"; d2 <= "0101"; d3 <= "0111"; d4 <= "0001"; -- 1756
    when "0000011011011101" => d1 <= "0111"; d2 <= "0101"; d3 <= "0111"; d4 <= "0001"; -- 1757
    when "0000011011011110" => d1 <= "1000"; d2 <= "0101"; d3 <= "0111"; d4 <= "0001"; -- 1758
    when "0000011011011111" => d1 <= "1001"; d2 <= "0101"; d3 <= "0111"; d4 <= "0001"; -- 1759
    when "0000011011100000" => d1 <= "0000"; d2 <= "0110"; d3 <= "0111"; d4 <= "0001"; -- 1760
    when "0000011011100001" => d1 <= "0001"; d2 <= "0110"; d3 <= "0111"; d4 <= "0001"; -- 1761
    when "0000011011100010" => d1 <= "0010"; d2 <= "0110"; d3 <= "0111"; d4 <= "0001"; -- 1762
    when "0000011011100011" => d1 <= "0011"; d2 <= "0110"; d3 <= "0111"; d4 <= "0001"; -- 1763
    when "0000011011100100" => d1 <= "0100"; d2 <= "0110"; d3 <= "0111"; d4 <= "0001"; -- 1764
    when "0000011011100101" => d1 <= "0101"; d2 <= "0110"; d3 <= "0111"; d4 <= "0001"; -- 1765
    when "0000011011100110" => d1 <= "0110"; d2 <= "0110"; d3 <= "0111"; d4 <= "0001"; -- 1766
    when "0000011011100111" => d1 <= "0111"; d2 <= "0110"; d3 <= "0111"; d4 <= "0001"; -- 1767
    when "0000011011101000" => d1 <= "1000"; d2 <= "0110"; d3 <= "0111"; d4 <= "0001"; -- 1768
    when "0000011011101001" => d1 <= "1001"; d2 <= "0110"; d3 <= "0111"; d4 <= "0001"; -- 1769
    when "0000011011101010" => d1 <= "0000"; d2 <= "0111"; d3 <= "0111"; d4 <= "0001"; -- 1770
    when "0000011011101011" => d1 <= "0001"; d2 <= "0111"; d3 <= "0111"; d4 <= "0001"; -- 1771
    when "0000011011101100" => d1 <= "0010"; d2 <= "0111"; d3 <= "0111"; d4 <= "0001"; -- 1772
    when "0000011011101101" => d1 <= "0011"; d2 <= "0111"; d3 <= "0111"; d4 <= "0001"; -- 1773
    when "0000011011101110" => d1 <= "0100"; d2 <= "0111"; d3 <= "0111"; d4 <= "0001"; -- 1774
    when "0000011011101111" => d1 <= "0101"; d2 <= "0111"; d3 <= "0111"; d4 <= "0001"; -- 1775
    when "0000011011110000" => d1 <= "0110"; d2 <= "0111"; d3 <= "0111"; d4 <= "0001"; -- 1776
    when "0000011011110001" => d1 <= "0111"; d2 <= "0111"; d3 <= "0111"; d4 <= "0001"; -- 1777
    when "0000011011110010" => d1 <= "1000"; d2 <= "0111"; d3 <= "0111"; d4 <= "0001"; -- 1778
    when "0000011011110011" => d1 <= "1001"; d2 <= "0111"; d3 <= "0111"; d4 <= "0001"; -- 1779
    when "0000011011110100" => d1 <= "0000"; d2 <= "1000"; d3 <= "0111"; d4 <= "0001"; -- 1780
    when "0000011011110101" => d1 <= "0001"; d2 <= "1000"; d3 <= "0111"; d4 <= "0001"; -- 1781
    when "0000011011110110" => d1 <= "0010"; d2 <= "1000"; d3 <= "0111"; d4 <= "0001"; -- 1782
    when "0000011011110111" => d1 <= "0011"; d2 <= "1000"; d3 <= "0111"; d4 <= "0001"; -- 1783
    when "0000011011111000" => d1 <= "0100"; d2 <= "1000"; d3 <= "0111"; d4 <= "0001"; -- 1784
    when "0000011011111001" => d1 <= "0101"; d2 <= "1000"; d3 <= "0111"; d4 <= "0001"; -- 1785
    when "0000011011111010" => d1 <= "0110"; d2 <= "1000"; d3 <= "0111"; d4 <= "0001"; -- 1786
    when "0000011011111011" => d1 <= "0111"; d2 <= "1000"; d3 <= "0111"; d4 <= "0001"; -- 1787
    when "0000011011111100" => d1 <= "1000"; d2 <= "1000"; d3 <= "0111"; d4 <= "0001"; -- 1788
    when "0000011011111101" => d1 <= "1001"; d2 <= "1000"; d3 <= "0111"; d4 <= "0001"; -- 1789
    when "0000011011111110" => d1 <= "0000"; d2 <= "1001"; d3 <= "0111"; d4 <= "0001"; -- 1790
    when "0000011011111111" => d1 <= "0001"; d2 <= "1001"; d3 <= "0111"; d4 <= "0001"; -- 1791
    when "0000011100000000" => d1 <= "0010"; d2 <= "1001"; d3 <= "0111"; d4 <= "0001"; -- 1792
    when "0000011100000001" => d1 <= "0011"; d2 <= "1001"; d3 <= "0111"; d4 <= "0001"; -- 1793
    when "0000011100000010" => d1 <= "0100"; d2 <= "1001"; d3 <= "0111"; d4 <= "0001"; -- 1794
    when "0000011100000011" => d1 <= "0101"; d2 <= "1001"; d3 <= "0111"; d4 <= "0001"; -- 1795
    when "0000011100000100" => d1 <= "0110"; d2 <= "1001"; d3 <= "0111"; d4 <= "0001"; -- 1796
    when "0000011100000101" => d1 <= "0111"; d2 <= "1001"; d3 <= "0111"; d4 <= "0001"; -- 1797
    when "0000011100000110" => d1 <= "1000"; d2 <= "1001"; d3 <= "0111"; d4 <= "0001"; -- 1798
    when "0000011100000111" => d1 <= "1001"; d2 <= "1001"; d3 <= "0111"; d4 <= "0001"; -- 1799
    when "0000011100001000" => d1 <= "0000"; d2 <= "0000"; d3 <= "1000"; d4 <= "0001"; -- 1800
    when "0000011100001001" => d1 <= "0001"; d2 <= "0000"; d3 <= "1000"; d4 <= "0001"; -- 1801
    when "0000011100001010" => d1 <= "0010"; d2 <= "0000"; d3 <= "1000"; d4 <= "0001"; -- 1802
    when "0000011100001011" => d1 <= "0011"; d2 <= "0000"; d3 <= "1000"; d4 <= "0001"; -- 1803
    when "0000011100001100" => d1 <= "0100"; d2 <= "0000"; d3 <= "1000"; d4 <= "0001"; -- 1804
    when "0000011100001101" => d1 <= "0101"; d2 <= "0000"; d3 <= "1000"; d4 <= "0001"; -- 1805
    when "0000011100001110" => d1 <= "0110"; d2 <= "0000"; d3 <= "1000"; d4 <= "0001"; -- 1806
    when "0000011100001111" => d1 <= "0111"; d2 <= "0000"; d3 <= "1000"; d4 <= "0001"; -- 1807
    when "0000011100010000" => d1 <= "1000"; d2 <= "0000"; d3 <= "1000"; d4 <= "0001"; -- 1808
    when "0000011100010001" => d1 <= "1001"; d2 <= "0000"; d3 <= "1000"; d4 <= "0001"; -- 1809
    when "0000011100010010" => d1 <= "0000"; d2 <= "0001"; d3 <= "1000"; d4 <= "0001"; -- 1810
    when "0000011100010011" => d1 <= "0001"; d2 <= "0001"; d3 <= "1000"; d4 <= "0001"; -- 1811
    when "0000011100010100" => d1 <= "0010"; d2 <= "0001"; d3 <= "1000"; d4 <= "0001"; -- 1812
    when "0000011100010101" => d1 <= "0011"; d2 <= "0001"; d3 <= "1000"; d4 <= "0001"; -- 1813
    when "0000011100010110" => d1 <= "0100"; d2 <= "0001"; d3 <= "1000"; d4 <= "0001"; -- 1814
    when "0000011100010111" => d1 <= "0101"; d2 <= "0001"; d3 <= "1000"; d4 <= "0001"; -- 1815
    when "0000011100011000" => d1 <= "0110"; d2 <= "0001"; d3 <= "1000"; d4 <= "0001"; -- 1816
    when "0000011100011001" => d1 <= "0111"; d2 <= "0001"; d3 <= "1000"; d4 <= "0001"; -- 1817
    when "0000011100011010" => d1 <= "1000"; d2 <= "0001"; d3 <= "1000"; d4 <= "0001"; -- 1818
    when "0000011100011011" => d1 <= "1001"; d2 <= "0001"; d3 <= "1000"; d4 <= "0001"; -- 1819
    when "0000011100011100" => d1 <= "0000"; d2 <= "0010"; d3 <= "1000"; d4 <= "0001"; -- 1820
    when "0000011100011101" => d1 <= "0001"; d2 <= "0010"; d3 <= "1000"; d4 <= "0001"; -- 1821
    when "0000011100011110" => d1 <= "0010"; d2 <= "0010"; d3 <= "1000"; d4 <= "0001"; -- 1822
    when "0000011100011111" => d1 <= "0011"; d2 <= "0010"; d3 <= "1000"; d4 <= "0001"; -- 1823
    when "0000011100100000" => d1 <= "0100"; d2 <= "0010"; d3 <= "1000"; d4 <= "0001"; -- 1824
    when "0000011100100001" => d1 <= "0101"; d2 <= "0010"; d3 <= "1000"; d4 <= "0001"; -- 1825
    when "0000011100100010" => d1 <= "0110"; d2 <= "0010"; d3 <= "1000"; d4 <= "0001"; -- 1826
    when "0000011100100011" => d1 <= "0111"; d2 <= "0010"; d3 <= "1000"; d4 <= "0001"; -- 1827
    when "0000011100100100" => d1 <= "1000"; d2 <= "0010"; d3 <= "1000"; d4 <= "0001"; -- 1828
    when "0000011100100101" => d1 <= "1001"; d2 <= "0010"; d3 <= "1000"; d4 <= "0001"; -- 1829
    when "0000011100100110" => d1 <= "0000"; d2 <= "0011"; d3 <= "1000"; d4 <= "0001"; -- 1830
    when "0000011100100111" => d1 <= "0001"; d2 <= "0011"; d3 <= "1000"; d4 <= "0001"; -- 1831
    when "0000011100101000" => d1 <= "0010"; d2 <= "0011"; d3 <= "1000"; d4 <= "0001"; -- 1832
    when "0000011100101001" => d1 <= "0011"; d2 <= "0011"; d3 <= "1000"; d4 <= "0001"; -- 1833
    when "0000011100101010" => d1 <= "0100"; d2 <= "0011"; d3 <= "1000"; d4 <= "0001"; -- 1834
    when "0000011100101011" => d1 <= "0101"; d2 <= "0011"; d3 <= "1000"; d4 <= "0001"; -- 1835
    when "0000011100101100" => d1 <= "0110"; d2 <= "0011"; d3 <= "1000"; d4 <= "0001"; -- 1836
    when "0000011100101101" => d1 <= "0111"; d2 <= "0011"; d3 <= "1000"; d4 <= "0001"; -- 1837
    when "0000011100101110" => d1 <= "1000"; d2 <= "0011"; d3 <= "1000"; d4 <= "0001"; -- 1838
    when "0000011100101111" => d1 <= "1001"; d2 <= "0011"; d3 <= "1000"; d4 <= "0001"; -- 1839
    when "0000011100110000" => d1 <= "0000"; d2 <= "0100"; d3 <= "1000"; d4 <= "0001"; -- 1840
    when "0000011100110001" => d1 <= "0001"; d2 <= "0100"; d3 <= "1000"; d4 <= "0001"; -- 1841
    when "0000011100110010" => d1 <= "0010"; d2 <= "0100"; d3 <= "1000"; d4 <= "0001"; -- 1842
    when "0000011100110011" => d1 <= "0011"; d2 <= "0100"; d3 <= "1000"; d4 <= "0001"; -- 1843
    when "0000011100110100" => d1 <= "0100"; d2 <= "0100"; d3 <= "1000"; d4 <= "0001"; -- 1844
    when "0000011100110101" => d1 <= "0101"; d2 <= "0100"; d3 <= "1000"; d4 <= "0001"; -- 1845
    when "0000011100110110" => d1 <= "0110"; d2 <= "0100"; d3 <= "1000"; d4 <= "0001"; -- 1846
    when "0000011100110111" => d1 <= "0111"; d2 <= "0100"; d3 <= "1000"; d4 <= "0001"; -- 1847
    when "0000011100111000" => d1 <= "1000"; d2 <= "0100"; d3 <= "1000"; d4 <= "0001"; -- 1848
    when "0000011100111001" => d1 <= "1001"; d2 <= "0100"; d3 <= "1000"; d4 <= "0001"; -- 1849
    when "0000011100111010" => d1 <= "0000"; d2 <= "0101"; d3 <= "1000"; d4 <= "0001"; -- 1850
    when "0000011100111011" => d1 <= "0001"; d2 <= "0101"; d3 <= "1000"; d4 <= "0001"; -- 1851
    when "0000011100111100" => d1 <= "0010"; d2 <= "0101"; d3 <= "1000"; d4 <= "0001"; -- 1852
    when "0000011100111101" => d1 <= "0011"; d2 <= "0101"; d3 <= "1000"; d4 <= "0001"; -- 1853
    when "0000011100111110" => d1 <= "0100"; d2 <= "0101"; d3 <= "1000"; d4 <= "0001"; -- 1854
    when "0000011100111111" => d1 <= "0101"; d2 <= "0101"; d3 <= "1000"; d4 <= "0001"; -- 1855
    when "0000011101000000" => d1 <= "0110"; d2 <= "0101"; d3 <= "1000"; d4 <= "0001"; -- 1856
    when "0000011101000001" => d1 <= "0111"; d2 <= "0101"; d3 <= "1000"; d4 <= "0001"; -- 1857
    when "0000011101000010" => d1 <= "1000"; d2 <= "0101"; d3 <= "1000"; d4 <= "0001"; -- 1858
    when "0000011101000011" => d1 <= "1001"; d2 <= "0101"; d3 <= "1000"; d4 <= "0001"; -- 1859
    when "0000011101000100" => d1 <= "0000"; d2 <= "0110"; d3 <= "1000"; d4 <= "0001"; -- 1860
    when "0000011101000101" => d1 <= "0001"; d2 <= "0110"; d3 <= "1000"; d4 <= "0001"; -- 1861
    when "0000011101000110" => d1 <= "0010"; d2 <= "0110"; d3 <= "1000"; d4 <= "0001"; -- 1862
    when "0000011101000111" => d1 <= "0011"; d2 <= "0110"; d3 <= "1000"; d4 <= "0001"; -- 1863
    when "0000011101001000" => d1 <= "0100"; d2 <= "0110"; d3 <= "1000"; d4 <= "0001"; -- 1864
    when "0000011101001001" => d1 <= "0101"; d2 <= "0110"; d3 <= "1000"; d4 <= "0001"; -- 1865
    when "0000011101001010" => d1 <= "0110"; d2 <= "0110"; d3 <= "1000"; d4 <= "0001"; -- 1866
    when "0000011101001011" => d1 <= "0111"; d2 <= "0110"; d3 <= "1000"; d4 <= "0001"; -- 1867
    when "0000011101001100" => d1 <= "1000"; d2 <= "0110"; d3 <= "1000"; d4 <= "0001"; -- 1868
    when "0000011101001101" => d1 <= "1001"; d2 <= "0110"; d3 <= "1000"; d4 <= "0001"; -- 1869
    when "0000011101001110" => d1 <= "0000"; d2 <= "0111"; d3 <= "1000"; d4 <= "0001"; -- 1870
    when "0000011101001111" => d1 <= "0001"; d2 <= "0111"; d3 <= "1000"; d4 <= "0001"; -- 1871
    when "0000011101010000" => d1 <= "0010"; d2 <= "0111"; d3 <= "1000"; d4 <= "0001"; -- 1872
    when "0000011101010001" => d1 <= "0011"; d2 <= "0111"; d3 <= "1000"; d4 <= "0001"; -- 1873
    when "0000011101010010" => d1 <= "0100"; d2 <= "0111"; d3 <= "1000"; d4 <= "0001"; -- 1874
    when "0000011101010011" => d1 <= "0101"; d2 <= "0111"; d3 <= "1000"; d4 <= "0001"; -- 1875
    when "0000011101010100" => d1 <= "0110"; d2 <= "0111"; d3 <= "1000"; d4 <= "0001"; -- 1876
    when "0000011101010101" => d1 <= "0111"; d2 <= "0111"; d3 <= "1000"; d4 <= "0001"; -- 1877
    when "0000011101010110" => d1 <= "1000"; d2 <= "0111"; d3 <= "1000"; d4 <= "0001"; -- 1878
    when "0000011101010111" => d1 <= "1001"; d2 <= "0111"; d3 <= "1000"; d4 <= "0001"; -- 1879
    when "0000011101011000" => d1 <= "0000"; d2 <= "1000"; d3 <= "1000"; d4 <= "0001"; -- 1880
    when "0000011101011001" => d1 <= "0001"; d2 <= "1000"; d3 <= "1000"; d4 <= "0001"; -- 1881
    when "0000011101011010" => d1 <= "0010"; d2 <= "1000"; d3 <= "1000"; d4 <= "0001"; -- 1882
    when "0000011101011011" => d1 <= "0011"; d2 <= "1000"; d3 <= "1000"; d4 <= "0001"; -- 1883
    when "0000011101011100" => d1 <= "0100"; d2 <= "1000"; d3 <= "1000"; d4 <= "0001"; -- 1884
    when "0000011101011101" => d1 <= "0101"; d2 <= "1000"; d3 <= "1000"; d4 <= "0001"; -- 1885
    when "0000011101011110" => d1 <= "0110"; d2 <= "1000"; d3 <= "1000"; d4 <= "0001"; -- 1886
    when "0000011101011111" => d1 <= "0111"; d2 <= "1000"; d3 <= "1000"; d4 <= "0001"; -- 1887
    when "0000011101100000" => d1 <= "1000"; d2 <= "1000"; d3 <= "1000"; d4 <= "0001"; -- 1888
    when "0000011101100001" => d1 <= "1001"; d2 <= "1000"; d3 <= "1000"; d4 <= "0001"; -- 1889
    when "0000011101100010" => d1 <= "0000"; d2 <= "1001"; d3 <= "1000"; d4 <= "0001"; -- 1890
    when "0000011101100011" => d1 <= "0001"; d2 <= "1001"; d3 <= "1000"; d4 <= "0001"; -- 1891
    when "0000011101100100" => d1 <= "0010"; d2 <= "1001"; d3 <= "1000"; d4 <= "0001"; -- 1892
    when "0000011101100101" => d1 <= "0011"; d2 <= "1001"; d3 <= "1000"; d4 <= "0001"; -- 1893
    when "0000011101100110" => d1 <= "0100"; d2 <= "1001"; d3 <= "1000"; d4 <= "0001"; -- 1894
    when "0000011101100111" => d1 <= "0101"; d2 <= "1001"; d3 <= "1000"; d4 <= "0001"; -- 1895
    when "0000011101101000" => d1 <= "0110"; d2 <= "1001"; d3 <= "1000"; d4 <= "0001"; -- 1896
    when "0000011101101001" => d1 <= "0111"; d2 <= "1001"; d3 <= "1000"; d4 <= "0001"; -- 1897
    when "0000011101101010" => d1 <= "1000"; d2 <= "1001"; d3 <= "1000"; d4 <= "0001"; -- 1898
    when "0000011101101011" => d1 <= "1001"; d2 <= "1001"; d3 <= "1000"; d4 <= "0001"; -- 1899
    when "0000011101101100" => d1 <= "0000"; d2 <= "0000"; d3 <= "1001"; d4 <= "0001"; -- 1900
    when "0000011101101101" => d1 <= "0001"; d2 <= "0000"; d3 <= "1001"; d4 <= "0001"; -- 1901
    when "0000011101101110" => d1 <= "0010"; d2 <= "0000"; d3 <= "1001"; d4 <= "0001"; -- 1902
    when "0000011101101111" => d1 <= "0011"; d2 <= "0000"; d3 <= "1001"; d4 <= "0001"; -- 1903
    when "0000011101110000" => d1 <= "0100"; d2 <= "0000"; d3 <= "1001"; d4 <= "0001"; -- 1904
    when "0000011101110001" => d1 <= "0101"; d2 <= "0000"; d3 <= "1001"; d4 <= "0001"; -- 1905
    when "0000011101110010" => d1 <= "0110"; d2 <= "0000"; d3 <= "1001"; d4 <= "0001"; -- 1906
    when "0000011101110011" => d1 <= "0111"; d2 <= "0000"; d3 <= "1001"; d4 <= "0001"; -- 1907
    when "0000011101110100" => d1 <= "1000"; d2 <= "0000"; d3 <= "1001"; d4 <= "0001"; -- 1908
    when "0000011101110101" => d1 <= "1001"; d2 <= "0000"; d3 <= "1001"; d4 <= "0001"; -- 1909
    when "0000011101110110" => d1 <= "0000"; d2 <= "0001"; d3 <= "1001"; d4 <= "0001"; -- 1910
    when "0000011101110111" => d1 <= "0001"; d2 <= "0001"; d3 <= "1001"; d4 <= "0001"; -- 1911
    when "0000011101111000" => d1 <= "0010"; d2 <= "0001"; d3 <= "1001"; d4 <= "0001"; -- 1912
    when "0000011101111001" => d1 <= "0011"; d2 <= "0001"; d3 <= "1001"; d4 <= "0001"; -- 1913
    when "0000011101111010" => d1 <= "0100"; d2 <= "0001"; d3 <= "1001"; d4 <= "0001"; -- 1914
    when "0000011101111011" => d1 <= "0101"; d2 <= "0001"; d3 <= "1001"; d4 <= "0001"; -- 1915
    when "0000011101111100" => d1 <= "0110"; d2 <= "0001"; d3 <= "1001"; d4 <= "0001"; -- 1916
    when "0000011101111101" => d1 <= "0111"; d2 <= "0001"; d3 <= "1001"; d4 <= "0001"; -- 1917
    when "0000011101111110" => d1 <= "1000"; d2 <= "0001"; d3 <= "1001"; d4 <= "0001"; -- 1918
    when "0000011101111111" => d1 <= "1001"; d2 <= "0001"; d3 <= "1001"; d4 <= "0001"; -- 1919
    when "0000011110000000" => d1 <= "0000"; d2 <= "0010"; d3 <= "1001"; d4 <= "0001"; -- 1920
    when "0000011110000001" => d1 <= "0001"; d2 <= "0010"; d3 <= "1001"; d4 <= "0001"; -- 1921
    when "0000011110000010" => d1 <= "0010"; d2 <= "0010"; d3 <= "1001"; d4 <= "0001"; -- 1922
    when "0000011110000011" => d1 <= "0011"; d2 <= "0010"; d3 <= "1001"; d4 <= "0001"; -- 1923
    when "0000011110000100" => d1 <= "0100"; d2 <= "0010"; d3 <= "1001"; d4 <= "0001"; -- 1924
    when "0000011110000101" => d1 <= "0101"; d2 <= "0010"; d3 <= "1001"; d4 <= "0001"; -- 1925
    when "0000011110000110" => d1 <= "0110"; d2 <= "0010"; d3 <= "1001"; d4 <= "0001"; -- 1926
    when "0000011110000111" => d1 <= "0111"; d2 <= "0010"; d3 <= "1001"; d4 <= "0001"; -- 1927
    when "0000011110001000" => d1 <= "1000"; d2 <= "0010"; d3 <= "1001"; d4 <= "0001"; -- 1928
    when "0000011110001001" => d1 <= "1001"; d2 <= "0010"; d3 <= "1001"; d4 <= "0001"; -- 1929
    when "0000011110001010" => d1 <= "0000"; d2 <= "0011"; d3 <= "1001"; d4 <= "0001"; -- 1930
    when "0000011110001011" => d1 <= "0001"; d2 <= "0011"; d3 <= "1001"; d4 <= "0001"; -- 1931
    when "0000011110001100" => d1 <= "0010"; d2 <= "0011"; d3 <= "1001"; d4 <= "0001"; -- 1932
    when "0000011110001101" => d1 <= "0011"; d2 <= "0011"; d3 <= "1001"; d4 <= "0001"; -- 1933
    when "0000011110001110" => d1 <= "0100"; d2 <= "0011"; d3 <= "1001"; d4 <= "0001"; -- 1934
    when "0000011110001111" => d1 <= "0101"; d2 <= "0011"; d3 <= "1001"; d4 <= "0001"; -- 1935
    when "0000011110010000" => d1 <= "0110"; d2 <= "0011"; d3 <= "1001"; d4 <= "0001"; -- 1936
    when "0000011110010001" => d1 <= "0111"; d2 <= "0011"; d3 <= "1001"; d4 <= "0001"; -- 1937
    when "0000011110010010" => d1 <= "1000"; d2 <= "0011"; d3 <= "1001"; d4 <= "0001"; -- 1938
    when "0000011110010011" => d1 <= "1001"; d2 <= "0011"; d3 <= "1001"; d4 <= "0001"; -- 1939
    when "0000011110010100" => d1 <= "0000"; d2 <= "0100"; d3 <= "1001"; d4 <= "0001"; -- 1940
    when "0000011110010101" => d1 <= "0001"; d2 <= "0100"; d3 <= "1001"; d4 <= "0001"; -- 1941
    when "0000011110010110" => d1 <= "0010"; d2 <= "0100"; d3 <= "1001"; d4 <= "0001"; -- 1942
    when "0000011110010111" => d1 <= "0011"; d2 <= "0100"; d3 <= "1001"; d4 <= "0001"; -- 1943
    when "0000011110011000" => d1 <= "0100"; d2 <= "0100"; d3 <= "1001"; d4 <= "0001"; -- 1944
    when "0000011110011001" => d1 <= "0101"; d2 <= "0100"; d3 <= "1001"; d4 <= "0001"; -- 1945
    when "0000011110011010" => d1 <= "0110"; d2 <= "0100"; d3 <= "1001"; d4 <= "0001"; -- 1946
    when "0000011110011011" => d1 <= "0111"; d2 <= "0100"; d3 <= "1001"; d4 <= "0001"; -- 1947
    when "0000011110011100" => d1 <= "1000"; d2 <= "0100"; d3 <= "1001"; d4 <= "0001"; -- 1948
    when "0000011110011101" => d1 <= "1001"; d2 <= "0100"; d3 <= "1001"; d4 <= "0001"; -- 1949
    when "0000011110011110" => d1 <= "0000"; d2 <= "0101"; d3 <= "1001"; d4 <= "0001"; -- 1950
    when "0000011110011111" => d1 <= "0001"; d2 <= "0101"; d3 <= "1001"; d4 <= "0001"; -- 1951
    when "0000011110100000" => d1 <= "0010"; d2 <= "0101"; d3 <= "1001"; d4 <= "0001"; -- 1952
    when "0000011110100001" => d1 <= "0011"; d2 <= "0101"; d3 <= "1001"; d4 <= "0001"; -- 1953
    when "0000011110100010" => d1 <= "0100"; d2 <= "0101"; d3 <= "1001"; d4 <= "0001"; -- 1954
    when "0000011110100011" => d1 <= "0101"; d2 <= "0101"; d3 <= "1001"; d4 <= "0001"; -- 1955
    when "0000011110100100" => d1 <= "0110"; d2 <= "0101"; d3 <= "1001"; d4 <= "0001"; -- 1956
    when "0000011110100101" => d1 <= "0111"; d2 <= "0101"; d3 <= "1001"; d4 <= "0001"; -- 1957
    when "0000011110100110" => d1 <= "1000"; d2 <= "0101"; d3 <= "1001"; d4 <= "0001"; -- 1958
    when "0000011110100111" => d1 <= "1001"; d2 <= "0101"; d3 <= "1001"; d4 <= "0001"; -- 1959
    when "0000011110101000" => d1 <= "0000"; d2 <= "0110"; d3 <= "1001"; d4 <= "0001"; -- 1960
    when "0000011110101001" => d1 <= "0001"; d2 <= "0110"; d3 <= "1001"; d4 <= "0001"; -- 1961
    when "0000011110101010" => d1 <= "0010"; d2 <= "0110"; d3 <= "1001"; d4 <= "0001"; -- 1962
    when "0000011110101011" => d1 <= "0011"; d2 <= "0110"; d3 <= "1001"; d4 <= "0001"; -- 1963
    when "0000011110101100" => d1 <= "0100"; d2 <= "0110"; d3 <= "1001"; d4 <= "0001"; -- 1964
    when "0000011110101101" => d1 <= "0101"; d2 <= "0110"; d3 <= "1001"; d4 <= "0001"; -- 1965
    when "0000011110101110" => d1 <= "0110"; d2 <= "0110"; d3 <= "1001"; d4 <= "0001"; -- 1966
    when "0000011110101111" => d1 <= "0111"; d2 <= "0110"; d3 <= "1001"; d4 <= "0001"; -- 1967
    when "0000011110110000" => d1 <= "1000"; d2 <= "0110"; d3 <= "1001"; d4 <= "0001"; -- 1968
    when "0000011110110001" => d1 <= "1001"; d2 <= "0110"; d3 <= "1001"; d4 <= "0001"; -- 1969
    when "0000011110110010" => d1 <= "0000"; d2 <= "0111"; d3 <= "1001"; d4 <= "0001"; -- 1970
    when "0000011110110011" => d1 <= "0001"; d2 <= "0111"; d3 <= "1001"; d4 <= "0001"; -- 1971
    when "0000011110110100" => d1 <= "0010"; d2 <= "0111"; d3 <= "1001"; d4 <= "0001"; -- 1972
    when "0000011110110101" => d1 <= "0011"; d2 <= "0111"; d3 <= "1001"; d4 <= "0001"; -- 1973
    when "0000011110110110" => d1 <= "0100"; d2 <= "0111"; d3 <= "1001"; d4 <= "0001"; -- 1974
    when "0000011110110111" => d1 <= "0101"; d2 <= "0111"; d3 <= "1001"; d4 <= "0001"; -- 1975
    when "0000011110111000" => d1 <= "0110"; d2 <= "0111"; d3 <= "1001"; d4 <= "0001"; -- 1976
    when "0000011110111001" => d1 <= "0111"; d2 <= "0111"; d3 <= "1001"; d4 <= "0001"; -- 1977
    when "0000011110111010" => d1 <= "1000"; d2 <= "0111"; d3 <= "1001"; d4 <= "0001"; -- 1978
    when "0000011110111011" => d1 <= "1001"; d2 <= "0111"; d3 <= "1001"; d4 <= "0001"; -- 1979
    when "0000011110111100" => d1 <= "0000"; d2 <= "1000"; d3 <= "1001"; d4 <= "0001"; -- 1980
    when "0000011110111101" => d1 <= "0001"; d2 <= "1000"; d3 <= "1001"; d4 <= "0001"; -- 1981
    when "0000011110111110" => d1 <= "0010"; d2 <= "1000"; d3 <= "1001"; d4 <= "0001"; -- 1982
    when "0000011110111111" => d1 <= "0011"; d2 <= "1000"; d3 <= "1001"; d4 <= "0001"; -- 1983
    when "0000011111000000" => d1 <= "0100"; d2 <= "1000"; d3 <= "1001"; d4 <= "0001"; -- 1984
    when "0000011111000001" => d1 <= "0101"; d2 <= "1000"; d3 <= "1001"; d4 <= "0001"; -- 1985
    when "0000011111000010" => d1 <= "0110"; d2 <= "1000"; d3 <= "1001"; d4 <= "0001"; -- 1986
    when "0000011111000011" => d1 <= "0111"; d2 <= "1000"; d3 <= "1001"; d4 <= "0001"; -- 1987
    when "0000011111000100" => d1 <= "1000"; d2 <= "1000"; d3 <= "1001"; d4 <= "0001"; -- 1988
    when "0000011111000101" => d1 <= "1001"; d2 <= "1000"; d3 <= "1001"; d4 <= "0001"; -- 1989
    when "0000011111000110" => d1 <= "0000"; d2 <= "1001"; d3 <= "1001"; d4 <= "0001"; -- 1990
    when "0000011111000111" => d1 <= "0001"; d2 <= "1001"; d3 <= "1001"; d4 <= "0001"; -- 1991
    when "0000011111001000" => d1 <= "0010"; d2 <= "1001"; d3 <= "1001"; d4 <= "0001"; -- 1992
    when "0000011111001001" => d1 <= "0011"; d2 <= "1001"; d3 <= "1001"; d4 <= "0001"; -- 1993
    when "0000011111001010" => d1 <= "0100"; d2 <= "1001"; d3 <= "1001"; d4 <= "0001"; -- 1994
    when "0000011111001011" => d1 <= "0101"; d2 <= "1001"; d3 <= "1001"; d4 <= "0001"; -- 1995
    when "0000011111001100" => d1 <= "0110"; d2 <= "1001"; d3 <= "1001"; d4 <= "0001"; -- 1996
    when "0000011111001101" => d1 <= "0111"; d2 <= "1001"; d3 <= "1001"; d4 <= "0001"; -- 1997
    when "0000011111001110" => d1 <= "1000"; d2 <= "1001"; d3 <= "1001"; d4 <= "0001"; -- 1998
    when "0000011111001111" => d1 <= "1001"; d2 <= "1001"; d3 <= "1001"; d4 <= "0001"; -- 1999
    when "0000011111010000" => d1 <= "0000"; d2 <= "0000"; d3 <= "0000"; d4 <= "0010"; -- 2000
    when "0000011111010001" => d1 <= "0001"; d2 <= "0000"; d3 <= "0000"; d4 <= "0010"; -- 2001
    when "0000011111010010" => d1 <= "0010"; d2 <= "0000"; d3 <= "0000"; d4 <= "0010"; -- 2002
    when "0000011111010011" => d1 <= "0011"; d2 <= "0000"; d3 <= "0000"; d4 <= "0010"; -- 2003
    when "0000011111010100" => d1 <= "0100"; d2 <= "0000"; d3 <= "0000"; d4 <= "0010"; -- 2004
    when "0000011111010101" => d1 <= "0101"; d2 <= "0000"; d3 <= "0000"; d4 <= "0010"; -- 2005
    when "0000011111010110" => d1 <= "0110"; d2 <= "0000"; d3 <= "0000"; d4 <= "0010"; -- 2006
    when "0000011111010111" => d1 <= "0111"; d2 <= "0000"; d3 <= "0000"; d4 <= "0010"; -- 2007
    when "0000011111011000" => d1 <= "1000"; d2 <= "0000"; d3 <= "0000"; d4 <= "0010"; -- 2008
    when "0000011111011001" => d1 <= "1001"; d2 <= "0000"; d3 <= "0000"; d4 <= "0010"; -- 2009
    when "0000011111011010" => d1 <= "0000"; d2 <= "0001"; d3 <= "0000"; d4 <= "0010"; -- 2010
    when "0000011111011011" => d1 <= "0001"; d2 <= "0001"; d3 <= "0000"; d4 <= "0010"; -- 2011
    when "0000011111011100" => d1 <= "0010"; d2 <= "0001"; d3 <= "0000"; d4 <= "0010"; -- 2012
    when "0000011111011101" => d1 <= "0011"; d2 <= "0001"; d3 <= "0000"; d4 <= "0010"; -- 2013
    when "0000011111011110" => d1 <= "0100"; d2 <= "0001"; d3 <= "0000"; d4 <= "0010"; -- 2014
    when "0000011111011111" => d1 <= "0101"; d2 <= "0001"; d3 <= "0000"; d4 <= "0010"; -- 2015
    when "0000011111100000" => d1 <= "0110"; d2 <= "0001"; d3 <= "0000"; d4 <= "0010"; -- 2016
    when "0000011111100001" => d1 <= "0111"; d2 <= "0001"; d3 <= "0000"; d4 <= "0010"; -- 2017
    when "0000011111100010" => d1 <= "1000"; d2 <= "0001"; d3 <= "0000"; d4 <= "0010"; -- 2018
    when "0000011111100011" => d1 <= "1001"; d2 <= "0001"; d3 <= "0000"; d4 <= "0010"; -- 2019
    when "0000011111100100" => d1 <= "0000"; d2 <= "0010"; d3 <= "0000"; d4 <= "0010"; -- 2020
    when "0000011111100101" => d1 <= "0001"; d2 <= "0010"; d3 <= "0000"; d4 <= "0010"; -- 2021
    when "0000011111100110" => d1 <= "0010"; d2 <= "0010"; d3 <= "0000"; d4 <= "0010"; -- 2022
    when "0000011111100111" => d1 <= "0011"; d2 <= "0010"; d3 <= "0000"; d4 <= "0010"; -- 2023
    when "0000011111101000" => d1 <= "0100"; d2 <= "0010"; d3 <= "0000"; d4 <= "0010"; -- 2024
    when "0000011111101001" => d1 <= "0101"; d2 <= "0010"; d3 <= "0000"; d4 <= "0010"; -- 2025
    when "0000011111101010" => d1 <= "0110"; d2 <= "0010"; d3 <= "0000"; d4 <= "0010"; -- 2026
    when "0000011111101011" => d1 <= "0111"; d2 <= "0010"; d3 <= "0000"; d4 <= "0010"; -- 2027
    when "0000011111101100" => d1 <= "1000"; d2 <= "0010"; d3 <= "0000"; d4 <= "0010"; -- 2028
    when "0000011111101101" => d1 <= "1001"; d2 <= "0010"; d3 <= "0000"; d4 <= "0010"; -- 2029
    when "0000011111101110" => d1 <= "0000"; d2 <= "0011"; d3 <= "0000"; d4 <= "0010"; -- 2030
    when "0000011111101111" => d1 <= "0001"; d2 <= "0011"; d3 <= "0000"; d4 <= "0010"; -- 2031
    when "0000011111110000" => d1 <= "0010"; d2 <= "0011"; d3 <= "0000"; d4 <= "0010"; -- 2032
    when "0000011111110001" => d1 <= "0011"; d2 <= "0011"; d3 <= "0000"; d4 <= "0010"; -- 2033
    when "0000011111110010" => d1 <= "0100"; d2 <= "0011"; d3 <= "0000"; d4 <= "0010"; -- 2034
    when "0000011111110011" => d1 <= "0101"; d2 <= "0011"; d3 <= "0000"; d4 <= "0010"; -- 2035
    when "0000011111110100" => d1 <= "0110"; d2 <= "0011"; d3 <= "0000"; d4 <= "0010"; -- 2036
    when "0000011111110101" => d1 <= "0111"; d2 <= "0011"; d3 <= "0000"; d4 <= "0010"; -- 2037
    when "0000011111110110" => d1 <= "1000"; d2 <= "0011"; d3 <= "0000"; d4 <= "0010"; -- 2038
    when "0000011111110111" => d1 <= "1001"; d2 <= "0011"; d3 <= "0000"; d4 <= "0010"; -- 2039
    when "0000011111111000" => d1 <= "0000"; d2 <= "0100"; d3 <= "0000"; d4 <= "0010"; -- 2040
    when "0000011111111001" => d1 <= "0001"; d2 <= "0100"; d3 <= "0000"; d4 <= "0010"; -- 2041
    when "0000011111111010" => d1 <= "0010"; d2 <= "0100"; d3 <= "0000"; d4 <= "0010"; -- 2042
    when "0000011111111011" => d1 <= "0011"; d2 <= "0100"; d3 <= "0000"; d4 <= "0010"; -- 2043
    when "0000011111111100" => d1 <= "0100"; d2 <= "0100"; d3 <= "0000"; d4 <= "0010"; -- 2044
    when "0000011111111101" => d1 <= "0101"; d2 <= "0100"; d3 <= "0000"; d4 <= "0010"; -- 2045
    when "0000011111111110" => d1 <= "0110"; d2 <= "0100"; d3 <= "0000"; d4 <= "0010"; -- 2046
    when "0000011111111111" => d1 <= "0111"; d2 <= "0100"; d3 <= "0000"; d4 <= "0010"; -- 2047
    when "0000100000000000" => d1 <= "1000"; d2 <= "0100"; d3 <= "0000"; d4 <= "0010"; -- 2048
    when "0000100000000001" => d1 <= "1001"; d2 <= "0100"; d3 <= "0000"; d4 <= "0010"; -- 2049
    when "0000100000000010" => d1 <= "0000"; d2 <= "0101"; d3 <= "0000"; d4 <= "0010"; -- 2050
    when "0000100000000011" => d1 <= "0001"; d2 <= "0101"; d3 <= "0000"; d4 <= "0010"; -- 2051
    when "0000100000000100" => d1 <= "0010"; d2 <= "0101"; d3 <= "0000"; d4 <= "0010"; -- 2052
    when "0000100000000101" => d1 <= "0011"; d2 <= "0101"; d3 <= "0000"; d4 <= "0010"; -- 2053
    when "0000100000000110" => d1 <= "0100"; d2 <= "0101"; d3 <= "0000"; d4 <= "0010"; -- 2054
    when "0000100000000111" => d1 <= "0101"; d2 <= "0101"; d3 <= "0000"; d4 <= "0010"; -- 2055
    when "0000100000001000" => d1 <= "0110"; d2 <= "0101"; d3 <= "0000"; d4 <= "0010"; -- 2056
    when "0000100000001001" => d1 <= "0111"; d2 <= "0101"; d3 <= "0000"; d4 <= "0010"; -- 2057
    when "0000100000001010" => d1 <= "1000"; d2 <= "0101"; d3 <= "0000"; d4 <= "0010"; -- 2058
    when "0000100000001011" => d1 <= "1001"; d2 <= "0101"; d3 <= "0000"; d4 <= "0010"; -- 2059
    when "0000100000001100" => d1 <= "0000"; d2 <= "0110"; d3 <= "0000"; d4 <= "0010"; -- 2060
    when "0000100000001101" => d1 <= "0001"; d2 <= "0110"; d3 <= "0000"; d4 <= "0010"; -- 2061
    when "0000100000001110" => d1 <= "0010"; d2 <= "0110"; d3 <= "0000"; d4 <= "0010"; -- 2062
    when "0000100000001111" => d1 <= "0011"; d2 <= "0110"; d3 <= "0000"; d4 <= "0010"; -- 2063
    when "0000100000010000" => d1 <= "0100"; d2 <= "0110"; d3 <= "0000"; d4 <= "0010"; -- 2064
    when "0000100000010001" => d1 <= "0101"; d2 <= "0110"; d3 <= "0000"; d4 <= "0010"; -- 2065
    when "0000100000010010" => d1 <= "0110"; d2 <= "0110"; d3 <= "0000"; d4 <= "0010"; -- 2066
    when "0000100000010011" => d1 <= "0111"; d2 <= "0110"; d3 <= "0000"; d4 <= "0010"; -- 2067
    when "0000100000010100" => d1 <= "1000"; d2 <= "0110"; d3 <= "0000"; d4 <= "0010"; -- 2068
    when "0000100000010101" => d1 <= "1001"; d2 <= "0110"; d3 <= "0000"; d4 <= "0010"; -- 2069
    when "0000100000010110" => d1 <= "0000"; d2 <= "0111"; d3 <= "0000"; d4 <= "0010"; -- 2070
    when "0000100000010111" => d1 <= "0001"; d2 <= "0111"; d3 <= "0000"; d4 <= "0010"; -- 2071
    when "0000100000011000" => d1 <= "0010"; d2 <= "0111"; d3 <= "0000"; d4 <= "0010"; -- 2072
    when "0000100000011001" => d1 <= "0011"; d2 <= "0111"; d3 <= "0000"; d4 <= "0010"; -- 2073
    when "0000100000011010" => d1 <= "0100"; d2 <= "0111"; d3 <= "0000"; d4 <= "0010"; -- 2074
    when "0000100000011011" => d1 <= "0101"; d2 <= "0111"; d3 <= "0000"; d4 <= "0010"; -- 2075
    when "0000100000011100" => d1 <= "0110"; d2 <= "0111"; d3 <= "0000"; d4 <= "0010"; -- 2076
    when "0000100000011101" => d1 <= "0111"; d2 <= "0111"; d3 <= "0000"; d4 <= "0010"; -- 2077
    when "0000100000011110" => d1 <= "1000"; d2 <= "0111"; d3 <= "0000"; d4 <= "0010"; -- 2078
    when "0000100000011111" => d1 <= "1001"; d2 <= "0111"; d3 <= "0000"; d4 <= "0010"; -- 2079
    when "0000100000100000" => d1 <= "0000"; d2 <= "1000"; d3 <= "0000"; d4 <= "0010"; -- 2080
    when "0000100000100001" => d1 <= "0001"; d2 <= "1000"; d3 <= "0000"; d4 <= "0010"; -- 2081
    when "0000100000100010" => d1 <= "0010"; d2 <= "1000"; d3 <= "0000"; d4 <= "0010"; -- 2082
    when "0000100000100011" => d1 <= "0011"; d2 <= "1000"; d3 <= "0000"; d4 <= "0010"; -- 2083
    when "0000100000100100" => d1 <= "0100"; d2 <= "1000"; d3 <= "0000"; d4 <= "0010"; -- 2084
    when "0000100000100101" => d1 <= "0101"; d2 <= "1000"; d3 <= "0000"; d4 <= "0010"; -- 2085
    when "0000100000100110" => d1 <= "0110"; d2 <= "1000"; d3 <= "0000"; d4 <= "0010"; -- 2086
    when "0000100000100111" => d1 <= "0111"; d2 <= "1000"; d3 <= "0000"; d4 <= "0010"; -- 2087
    when "0000100000101000" => d1 <= "1000"; d2 <= "1000"; d3 <= "0000"; d4 <= "0010"; -- 2088
    when "0000100000101001" => d1 <= "1001"; d2 <= "1000"; d3 <= "0000"; d4 <= "0010"; -- 2089
    when "0000100000101010" => d1 <= "0000"; d2 <= "1001"; d3 <= "0000"; d4 <= "0010"; -- 2090
    when "0000100000101011" => d1 <= "0001"; d2 <= "1001"; d3 <= "0000"; d4 <= "0010"; -- 2091
    when "0000100000101100" => d1 <= "0010"; d2 <= "1001"; d3 <= "0000"; d4 <= "0010"; -- 2092
    when "0000100000101101" => d1 <= "0011"; d2 <= "1001"; d3 <= "0000"; d4 <= "0010"; -- 2093
    when "0000100000101110" => d1 <= "0100"; d2 <= "1001"; d3 <= "0000"; d4 <= "0010"; -- 2094
    when "0000100000101111" => d1 <= "0101"; d2 <= "1001"; d3 <= "0000"; d4 <= "0010"; -- 2095
    when "0000100000110000" => d1 <= "0110"; d2 <= "1001"; d3 <= "0000"; d4 <= "0010"; -- 2096
    when "0000100000110001" => d1 <= "0111"; d2 <= "1001"; d3 <= "0000"; d4 <= "0010"; -- 2097
    when "0000100000110010" => d1 <= "1000"; d2 <= "1001"; d3 <= "0000"; d4 <= "0010"; -- 2098
    when "0000100000110011" => d1 <= "1001"; d2 <= "1001"; d3 <= "0000"; d4 <= "0010"; -- 2099
    when "0000100000110100" => d1 <= "0000"; d2 <= "0000"; d3 <= "0001"; d4 <= "0010"; -- 2100
    when "0000100000110101" => d1 <= "0001"; d2 <= "0000"; d3 <= "0001"; d4 <= "0010"; -- 2101
    when "0000100000110110" => d1 <= "0010"; d2 <= "0000"; d3 <= "0001"; d4 <= "0010"; -- 2102
    when "0000100000110111" => d1 <= "0011"; d2 <= "0000"; d3 <= "0001"; d4 <= "0010"; -- 2103
    when "0000100000111000" => d1 <= "0100"; d2 <= "0000"; d3 <= "0001"; d4 <= "0010"; -- 2104
    when "0000100000111001" => d1 <= "0101"; d2 <= "0000"; d3 <= "0001"; d4 <= "0010"; -- 2105
    when "0000100000111010" => d1 <= "0110"; d2 <= "0000"; d3 <= "0001"; d4 <= "0010"; -- 2106
    when "0000100000111011" => d1 <= "0111"; d2 <= "0000"; d3 <= "0001"; d4 <= "0010"; -- 2107
    when "0000100000111100" => d1 <= "1000"; d2 <= "0000"; d3 <= "0001"; d4 <= "0010"; -- 2108
    when "0000100000111101" => d1 <= "1001"; d2 <= "0000"; d3 <= "0001"; d4 <= "0010"; -- 2109
    when "0000100000111110" => d1 <= "0000"; d2 <= "0001"; d3 <= "0001"; d4 <= "0010"; -- 2110
    when "0000100000111111" => d1 <= "0001"; d2 <= "0001"; d3 <= "0001"; d4 <= "0010"; -- 2111
    when "0000100001000000" => d1 <= "0010"; d2 <= "0001"; d3 <= "0001"; d4 <= "0010"; -- 2112
    when "0000100001000001" => d1 <= "0011"; d2 <= "0001"; d3 <= "0001"; d4 <= "0010"; -- 2113
    when "0000100001000010" => d1 <= "0100"; d2 <= "0001"; d3 <= "0001"; d4 <= "0010"; -- 2114
    when "0000100001000011" => d1 <= "0101"; d2 <= "0001"; d3 <= "0001"; d4 <= "0010"; -- 2115
    when "0000100001000100" => d1 <= "0110"; d2 <= "0001"; d3 <= "0001"; d4 <= "0010"; -- 2116
    when "0000100001000101" => d1 <= "0111"; d2 <= "0001"; d3 <= "0001"; d4 <= "0010"; -- 2117
    when "0000100001000110" => d1 <= "1000"; d2 <= "0001"; d3 <= "0001"; d4 <= "0010"; -- 2118
    when "0000100001000111" => d1 <= "1001"; d2 <= "0001"; d3 <= "0001"; d4 <= "0010"; -- 2119
    when "0000100001001000" => d1 <= "0000"; d2 <= "0010"; d3 <= "0001"; d4 <= "0010"; -- 2120
    when "0000100001001001" => d1 <= "0001"; d2 <= "0010"; d3 <= "0001"; d4 <= "0010"; -- 2121
    when "0000100001001010" => d1 <= "0010"; d2 <= "0010"; d3 <= "0001"; d4 <= "0010"; -- 2122
    when "0000100001001011" => d1 <= "0011"; d2 <= "0010"; d3 <= "0001"; d4 <= "0010"; -- 2123
    when "0000100001001100" => d1 <= "0100"; d2 <= "0010"; d3 <= "0001"; d4 <= "0010"; -- 2124
    when "0000100001001101" => d1 <= "0101"; d2 <= "0010"; d3 <= "0001"; d4 <= "0010"; -- 2125
    when "0000100001001110" => d1 <= "0110"; d2 <= "0010"; d3 <= "0001"; d4 <= "0010"; -- 2126
    when "0000100001001111" => d1 <= "0111"; d2 <= "0010"; d3 <= "0001"; d4 <= "0010"; -- 2127
    when "0000100001010000" => d1 <= "1000"; d2 <= "0010"; d3 <= "0001"; d4 <= "0010"; -- 2128
    when "0000100001010001" => d1 <= "1001"; d2 <= "0010"; d3 <= "0001"; d4 <= "0010"; -- 2129
    when "0000100001010010" => d1 <= "0000"; d2 <= "0011"; d3 <= "0001"; d4 <= "0010"; -- 2130
    when "0000100001010011" => d1 <= "0001"; d2 <= "0011"; d3 <= "0001"; d4 <= "0010"; -- 2131
    when "0000100001010100" => d1 <= "0010"; d2 <= "0011"; d3 <= "0001"; d4 <= "0010"; -- 2132
    when "0000100001010101" => d1 <= "0011"; d2 <= "0011"; d3 <= "0001"; d4 <= "0010"; -- 2133
    when "0000100001010110" => d1 <= "0100"; d2 <= "0011"; d3 <= "0001"; d4 <= "0010"; -- 2134
    when "0000100001010111" => d1 <= "0101"; d2 <= "0011"; d3 <= "0001"; d4 <= "0010"; -- 2135
    when "0000100001011000" => d1 <= "0110"; d2 <= "0011"; d3 <= "0001"; d4 <= "0010"; -- 2136
    when "0000100001011001" => d1 <= "0111"; d2 <= "0011"; d3 <= "0001"; d4 <= "0010"; -- 2137
    when "0000100001011010" => d1 <= "1000"; d2 <= "0011"; d3 <= "0001"; d4 <= "0010"; -- 2138
    when "0000100001011011" => d1 <= "1001"; d2 <= "0011"; d3 <= "0001"; d4 <= "0010"; -- 2139
    when "0000100001011100" => d1 <= "0000"; d2 <= "0100"; d3 <= "0001"; d4 <= "0010"; -- 2140
    when "0000100001011101" => d1 <= "0001"; d2 <= "0100"; d3 <= "0001"; d4 <= "0010"; -- 2141
    when "0000100001011110" => d1 <= "0010"; d2 <= "0100"; d3 <= "0001"; d4 <= "0010"; -- 2142
    when "0000100001011111" => d1 <= "0011"; d2 <= "0100"; d3 <= "0001"; d4 <= "0010"; -- 2143
    when "0000100001100000" => d1 <= "0100"; d2 <= "0100"; d3 <= "0001"; d4 <= "0010"; -- 2144
    when "0000100001100001" => d1 <= "0101"; d2 <= "0100"; d3 <= "0001"; d4 <= "0010"; -- 2145
    when "0000100001100010" => d1 <= "0110"; d2 <= "0100"; d3 <= "0001"; d4 <= "0010"; -- 2146
    when "0000100001100011" => d1 <= "0111"; d2 <= "0100"; d3 <= "0001"; d4 <= "0010"; -- 2147
    when "0000100001100100" => d1 <= "1000"; d2 <= "0100"; d3 <= "0001"; d4 <= "0010"; -- 2148
    when "0000100001100101" => d1 <= "1001"; d2 <= "0100"; d3 <= "0001"; d4 <= "0010"; -- 2149
    when "0000100001100110" => d1 <= "0000"; d2 <= "0101"; d3 <= "0001"; d4 <= "0010"; -- 2150
    when "0000100001100111" => d1 <= "0001"; d2 <= "0101"; d3 <= "0001"; d4 <= "0010"; -- 2151
    when "0000100001101000" => d1 <= "0010"; d2 <= "0101"; d3 <= "0001"; d4 <= "0010"; -- 2152
    when "0000100001101001" => d1 <= "0011"; d2 <= "0101"; d3 <= "0001"; d4 <= "0010"; -- 2153
    when "0000100001101010" => d1 <= "0100"; d2 <= "0101"; d3 <= "0001"; d4 <= "0010"; -- 2154
    when "0000100001101011" => d1 <= "0101"; d2 <= "0101"; d3 <= "0001"; d4 <= "0010"; -- 2155
    when "0000100001101100" => d1 <= "0110"; d2 <= "0101"; d3 <= "0001"; d4 <= "0010"; -- 2156
    when "0000100001101101" => d1 <= "0111"; d2 <= "0101"; d3 <= "0001"; d4 <= "0010"; -- 2157
    when "0000100001101110" => d1 <= "1000"; d2 <= "0101"; d3 <= "0001"; d4 <= "0010"; -- 2158
    when "0000100001101111" => d1 <= "1001"; d2 <= "0101"; d3 <= "0001"; d4 <= "0010"; -- 2159
    when "0000100001110000" => d1 <= "0000"; d2 <= "0110"; d3 <= "0001"; d4 <= "0010"; -- 2160
    when "0000100001110001" => d1 <= "0001"; d2 <= "0110"; d3 <= "0001"; d4 <= "0010"; -- 2161
    when "0000100001110010" => d1 <= "0010"; d2 <= "0110"; d3 <= "0001"; d4 <= "0010"; -- 2162
    when "0000100001110011" => d1 <= "0011"; d2 <= "0110"; d3 <= "0001"; d4 <= "0010"; -- 2163
    when "0000100001110100" => d1 <= "0100"; d2 <= "0110"; d3 <= "0001"; d4 <= "0010"; -- 2164
    when "0000100001110101" => d1 <= "0101"; d2 <= "0110"; d3 <= "0001"; d4 <= "0010"; -- 2165
    when "0000100001110110" => d1 <= "0110"; d2 <= "0110"; d3 <= "0001"; d4 <= "0010"; -- 2166
    when "0000100001110111" => d1 <= "0111"; d2 <= "0110"; d3 <= "0001"; d4 <= "0010"; -- 2167
    when "0000100001111000" => d1 <= "1000"; d2 <= "0110"; d3 <= "0001"; d4 <= "0010"; -- 2168
    when "0000100001111001" => d1 <= "1001"; d2 <= "0110"; d3 <= "0001"; d4 <= "0010"; -- 2169
    when "0000100001111010" => d1 <= "0000"; d2 <= "0111"; d3 <= "0001"; d4 <= "0010"; -- 2170
    when "0000100001111011" => d1 <= "0001"; d2 <= "0111"; d3 <= "0001"; d4 <= "0010"; -- 2171
    when "0000100001111100" => d1 <= "0010"; d2 <= "0111"; d3 <= "0001"; d4 <= "0010"; -- 2172
    when "0000100001111101" => d1 <= "0011"; d2 <= "0111"; d3 <= "0001"; d4 <= "0010"; -- 2173
    when "0000100001111110" => d1 <= "0100"; d2 <= "0111"; d3 <= "0001"; d4 <= "0010"; -- 2174
    when "0000100001111111" => d1 <= "0101"; d2 <= "0111"; d3 <= "0001"; d4 <= "0010"; -- 2175
    when "0000100010000000" => d1 <= "0110"; d2 <= "0111"; d3 <= "0001"; d4 <= "0010"; -- 2176
    when "0000100010000001" => d1 <= "0111"; d2 <= "0111"; d3 <= "0001"; d4 <= "0010"; -- 2177
    when "0000100010000010" => d1 <= "1000"; d2 <= "0111"; d3 <= "0001"; d4 <= "0010"; -- 2178
    when "0000100010000011" => d1 <= "1001"; d2 <= "0111"; d3 <= "0001"; d4 <= "0010"; -- 2179
    when "0000100010000100" => d1 <= "0000"; d2 <= "1000"; d3 <= "0001"; d4 <= "0010"; -- 2180
    when "0000100010000101" => d1 <= "0001"; d2 <= "1000"; d3 <= "0001"; d4 <= "0010"; -- 2181
    when "0000100010000110" => d1 <= "0010"; d2 <= "1000"; d3 <= "0001"; d4 <= "0010"; -- 2182
    when "0000100010000111" => d1 <= "0011"; d2 <= "1000"; d3 <= "0001"; d4 <= "0010"; -- 2183
    when "0000100010001000" => d1 <= "0100"; d2 <= "1000"; d3 <= "0001"; d4 <= "0010"; -- 2184
    when "0000100010001001" => d1 <= "0101"; d2 <= "1000"; d3 <= "0001"; d4 <= "0010"; -- 2185
    when "0000100010001010" => d1 <= "0110"; d2 <= "1000"; d3 <= "0001"; d4 <= "0010"; -- 2186
    when "0000100010001011" => d1 <= "0111"; d2 <= "1000"; d3 <= "0001"; d4 <= "0010"; -- 2187
    when "0000100010001100" => d1 <= "1000"; d2 <= "1000"; d3 <= "0001"; d4 <= "0010"; -- 2188
    when "0000100010001101" => d1 <= "1001"; d2 <= "1000"; d3 <= "0001"; d4 <= "0010"; -- 2189
    when "0000100010001110" => d1 <= "0000"; d2 <= "1001"; d3 <= "0001"; d4 <= "0010"; -- 2190
    when "0000100010001111" => d1 <= "0001"; d2 <= "1001"; d3 <= "0001"; d4 <= "0010"; -- 2191
    when "0000100010010000" => d1 <= "0010"; d2 <= "1001"; d3 <= "0001"; d4 <= "0010"; -- 2192
    when "0000100010010001" => d1 <= "0011"; d2 <= "1001"; d3 <= "0001"; d4 <= "0010"; -- 2193
    when "0000100010010010" => d1 <= "0100"; d2 <= "1001"; d3 <= "0001"; d4 <= "0010"; -- 2194
    when "0000100010010011" => d1 <= "0101"; d2 <= "1001"; d3 <= "0001"; d4 <= "0010"; -- 2195
    when "0000100010010100" => d1 <= "0110"; d2 <= "1001"; d3 <= "0001"; d4 <= "0010"; -- 2196
    when "0000100010010101" => d1 <= "0111"; d2 <= "1001"; d3 <= "0001"; d4 <= "0010"; -- 2197
    when "0000100010010110" => d1 <= "1000"; d2 <= "1001"; d3 <= "0001"; d4 <= "0010"; -- 2198
    when "0000100010010111" => d1 <= "1001"; d2 <= "1001"; d3 <= "0001"; d4 <= "0010"; -- 2199
    when "0000100010011000" => d1 <= "0000"; d2 <= "0000"; d3 <= "0010"; d4 <= "0010"; -- 2200
    when "0000100010011001" => d1 <= "0001"; d2 <= "0000"; d3 <= "0010"; d4 <= "0010"; -- 2201
    when "0000100010011010" => d1 <= "0010"; d2 <= "0000"; d3 <= "0010"; d4 <= "0010"; -- 2202
    when "0000100010011011" => d1 <= "0011"; d2 <= "0000"; d3 <= "0010"; d4 <= "0010"; -- 2203
    when "0000100010011100" => d1 <= "0100"; d2 <= "0000"; d3 <= "0010"; d4 <= "0010"; -- 2204
    when "0000100010011101" => d1 <= "0101"; d2 <= "0000"; d3 <= "0010"; d4 <= "0010"; -- 2205
    when "0000100010011110" => d1 <= "0110"; d2 <= "0000"; d3 <= "0010"; d4 <= "0010"; -- 2206
    when "0000100010011111" => d1 <= "0111"; d2 <= "0000"; d3 <= "0010"; d4 <= "0010"; -- 2207
    when "0000100010100000" => d1 <= "1000"; d2 <= "0000"; d3 <= "0010"; d4 <= "0010"; -- 2208
    when "0000100010100001" => d1 <= "1001"; d2 <= "0000"; d3 <= "0010"; d4 <= "0010"; -- 2209
    when "0000100010100010" => d1 <= "0000"; d2 <= "0001"; d3 <= "0010"; d4 <= "0010"; -- 2210
    when "0000100010100011" => d1 <= "0001"; d2 <= "0001"; d3 <= "0010"; d4 <= "0010"; -- 2211
    when "0000100010100100" => d1 <= "0010"; d2 <= "0001"; d3 <= "0010"; d4 <= "0010"; -- 2212
    when "0000100010100101" => d1 <= "0011"; d2 <= "0001"; d3 <= "0010"; d4 <= "0010"; -- 2213
    when "0000100010100110" => d1 <= "0100"; d2 <= "0001"; d3 <= "0010"; d4 <= "0010"; -- 2214
    when "0000100010100111" => d1 <= "0101"; d2 <= "0001"; d3 <= "0010"; d4 <= "0010"; -- 2215
    when "0000100010101000" => d1 <= "0110"; d2 <= "0001"; d3 <= "0010"; d4 <= "0010"; -- 2216
    when "0000100010101001" => d1 <= "0111"; d2 <= "0001"; d3 <= "0010"; d4 <= "0010"; -- 2217
    when "0000100010101010" => d1 <= "1000"; d2 <= "0001"; d3 <= "0010"; d4 <= "0010"; -- 2218
    when "0000100010101011" => d1 <= "1001"; d2 <= "0001"; d3 <= "0010"; d4 <= "0010"; -- 2219
    when "0000100010101100" => d1 <= "0000"; d2 <= "0010"; d3 <= "0010"; d4 <= "0010"; -- 2220
    when "0000100010101101" => d1 <= "0001"; d2 <= "0010"; d3 <= "0010"; d4 <= "0010"; -- 2221
    when "0000100010101110" => d1 <= "0010"; d2 <= "0010"; d3 <= "0010"; d4 <= "0010"; -- 2222
    when "0000100010101111" => d1 <= "0011"; d2 <= "0010"; d3 <= "0010"; d4 <= "0010"; -- 2223
    when "0000100010110000" => d1 <= "0100"; d2 <= "0010"; d3 <= "0010"; d4 <= "0010"; -- 2224
    when "0000100010110001" => d1 <= "0101"; d2 <= "0010"; d3 <= "0010"; d4 <= "0010"; -- 2225
    when "0000100010110010" => d1 <= "0110"; d2 <= "0010"; d3 <= "0010"; d4 <= "0010"; -- 2226
    when "0000100010110011" => d1 <= "0111"; d2 <= "0010"; d3 <= "0010"; d4 <= "0010"; -- 2227
    when "0000100010110100" => d1 <= "1000"; d2 <= "0010"; d3 <= "0010"; d4 <= "0010"; -- 2228
    when "0000100010110101" => d1 <= "1001"; d2 <= "0010"; d3 <= "0010"; d4 <= "0010"; -- 2229
    when "0000100010110110" => d1 <= "0000"; d2 <= "0011"; d3 <= "0010"; d4 <= "0010"; -- 2230
    when "0000100010110111" => d1 <= "0001"; d2 <= "0011"; d3 <= "0010"; d4 <= "0010"; -- 2231
    when "0000100010111000" => d1 <= "0010"; d2 <= "0011"; d3 <= "0010"; d4 <= "0010"; -- 2232
    when "0000100010111001" => d1 <= "0011"; d2 <= "0011"; d3 <= "0010"; d4 <= "0010"; -- 2233
    when "0000100010111010" => d1 <= "0100"; d2 <= "0011"; d3 <= "0010"; d4 <= "0010"; -- 2234
    when "0000100010111011" => d1 <= "0101"; d2 <= "0011"; d3 <= "0010"; d4 <= "0010"; -- 2235
    when "0000100010111100" => d1 <= "0110"; d2 <= "0011"; d3 <= "0010"; d4 <= "0010"; -- 2236
    when "0000100010111101" => d1 <= "0111"; d2 <= "0011"; d3 <= "0010"; d4 <= "0010"; -- 2237
    when "0000100010111110" => d1 <= "1000"; d2 <= "0011"; d3 <= "0010"; d4 <= "0010"; -- 2238
    when "0000100010111111" => d1 <= "1001"; d2 <= "0011"; d3 <= "0010"; d4 <= "0010"; -- 2239
    when "0000100011000000" => d1 <= "0000"; d2 <= "0100"; d3 <= "0010"; d4 <= "0010"; -- 2240
    when "0000100011000001" => d1 <= "0001"; d2 <= "0100"; d3 <= "0010"; d4 <= "0010"; -- 2241
    when "0000100011000010" => d1 <= "0010"; d2 <= "0100"; d3 <= "0010"; d4 <= "0010"; -- 2242
    when "0000100011000011" => d1 <= "0011"; d2 <= "0100"; d3 <= "0010"; d4 <= "0010"; -- 2243
    when "0000100011000100" => d1 <= "0100"; d2 <= "0100"; d3 <= "0010"; d4 <= "0010"; -- 2244
    when "0000100011000101" => d1 <= "0101"; d2 <= "0100"; d3 <= "0010"; d4 <= "0010"; -- 2245
    when "0000100011000110" => d1 <= "0110"; d2 <= "0100"; d3 <= "0010"; d4 <= "0010"; -- 2246
    when "0000100011000111" => d1 <= "0111"; d2 <= "0100"; d3 <= "0010"; d4 <= "0010"; -- 2247
    when "0000100011001000" => d1 <= "1000"; d2 <= "0100"; d3 <= "0010"; d4 <= "0010"; -- 2248
    when "0000100011001001" => d1 <= "1001"; d2 <= "0100"; d3 <= "0010"; d4 <= "0010"; -- 2249
    when "0000100011001010" => d1 <= "0000"; d2 <= "0101"; d3 <= "0010"; d4 <= "0010"; -- 2250
    when "0000100011001011" => d1 <= "0001"; d2 <= "0101"; d3 <= "0010"; d4 <= "0010"; -- 2251
    when "0000100011001100" => d1 <= "0010"; d2 <= "0101"; d3 <= "0010"; d4 <= "0010"; -- 2252
    when "0000100011001101" => d1 <= "0011"; d2 <= "0101"; d3 <= "0010"; d4 <= "0010"; -- 2253
    when "0000100011001110" => d1 <= "0100"; d2 <= "0101"; d3 <= "0010"; d4 <= "0010"; -- 2254
    when "0000100011001111" => d1 <= "0101"; d2 <= "0101"; d3 <= "0010"; d4 <= "0010"; -- 2255
    when "0000100011010000" => d1 <= "0110"; d2 <= "0101"; d3 <= "0010"; d4 <= "0010"; -- 2256
    when "0000100011010001" => d1 <= "0111"; d2 <= "0101"; d3 <= "0010"; d4 <= "0010"; -- 2257
    when "0000100011010010" => d1 <= "1000"; d2 <= "0101"; d3 <= "0010"; d4 <= "0010"; -- 2258
    when "0000100011010011" => d1 <= "1001"; d2 <= "0101"; d3 <= "0010"; d4 <= "0010"; -- 2259
    when "0000100011010100" => d1 <= "0000"; d2 <= "0110"; d3 <= "0010"; d4 <= "0010"; -- 2260
    when "0000100011010101" => d1 <= "0001"; d2 <= "0110"; d3 <= "0010"; d4 <= "0010"; -- 2261
    when "0000100011010110" => d1 <= "0010"; d2 <= "0110"; d3 <= "0010"; d4 <= "0010"; -- 2262
    when "0000100011010111" => d1 <= "0011"; d2 <= "0110"; d3 <= "0010"; d4 <= "0010"; -- 2263
    when "0000100011011000" => d1 <= "0100"; d2 <= "0110"; d3 <= "0010"; d4 <= "0010"; -- 2264
    when "0000100011011001" => d1 <= "0101"; d2 <= "0110"; d3 <= "0010"; d4 <= "0010"; -- 2265
    when "0000100011011010" => d1 <= "0110"; d2 <= "0110"; d3 <= "0010"; d4 <= "0010"; -- 2266
    when "0000100011011011" => d1 <= "0111"; d2 <= "0110"; d3 <= "0010"; d4 <= "0010"; -- 2267
    when "0000100011011100" => d1 <= "1000"; d2 <= "0110"; d3 <= "0010"; d4 <= "0010"; -- 2268
    when "0000100011011101" => d1 <= "1001"; d2 <= "0110"; d3 <= "0010"; d4 <= "0010"; -- 2269
    when "0000100011011110" => d1 <= "0000"; d2 <= "0111"; d3 <= "0010"; d4 <= "0010"; -- 2270
    when "0000100011011111" => d1 <= "0001"; d2 <= "0111"; d3 <= "0010"; d4 <= "0010"; -- 2271
    when "0000100011100000" => d1 <= "0010"; d2 <= "0111"; d3 <= "0010"; d4 <= "0010"; -- 2272
    when "0000100011100001" => d1 <= "0011"; d2 <= "0111"; d3 <= "0010"; d4 <= "0010"; -- 2273
    when "0000100011100010" => d1 <= "0100"; d2 <= "0111"; d3 <= "0010"; d4 <= "0010"; -- 2274
    when "0000100011100011" => d1 <= "0101"; d2 <= "0111"; d3 <= "0010"; d4 <= "0010"; -- 2275
    when "0000100011100100" => d1 <= "0110"; d2 <= "0111"; d3 <= "0010"; d4 <= "0010"; -- 2276
    when "0000100011100101" => d1 <= "0111"; d2 <= "0111"; d3 <= "0010"; d4 <= "0010"; -- 2277
    when "0000100011100110" => d1 <= "1000"; d2 <= "0111"; d3 <= "0010"; d4 <= "0010"; -- 2278
    when "0000100011100111" => d1 <= "1001"; d2 <= "0111"; d3 <= "0010"; d4 <= "0010"; -- 2279
    when "0000100011101000" => d1 <= "0000"; d2 <= "1000"; d3 <= "0010"; d4 <= "0010"; -- 2280
    when "0000100011101001" => d1 <= "0001"; d2 <= "1000"; d3 <= "0010"; d4 <= "0010"; -- 2281
    when "0000100011101010" => d1 <= "0010"; d2 <= "1000"; d3 <= "0010"; d4 <= "0010"; -- 2282
    when "0000100011101011" => d1 <= "0011"; d2 <= "1000"; d3 <= "0010"; d4 <= "0010"; -- 2283
    when "0000100011101100" => d1 <= "0100"; d2 <= "1000"; d3 <= "0010"; d4 <= "0010"; -- 2284
    when "0000100011101101" => d1 <= "0101"; d2 <= "1000"; d3 <= "0010"; d4 <= "0010"; -- 2285
    when "0000100011101110" => d1 <= "0110"; d2 <= "1000"; d3 <= "0010"; d4 <= "0010"; -- 2286
    when "0000100011101111" => d1 <= "0111"; d2 <= "1000"; d3 <= "0010"; d4 <= "0010"; -- 2287
    when "0000100011110000" => d1 <= "1000"; d2 <= "1000"; d3 <= "0010"; d4 <= "0010"; -- 2288
    when "0000100011110001" => d1 <= "1001"; d2 <= "1000"; d3 <= "0010"; d4 <= "0010"; -- 2289
    when "0000100011110010" => d1 <= "0000"; d2 <= "1001"; d3 <= "0010"; d4 <= "0010"; -- 2290
    when "0000100011110011" => d1 <= "0001"; d2 <= "1001"; d3 <= "0010"; d4 <= "0010"; -- 2291
    when "0000100011110100" => d1 <= "0010"; d2 <= "1001"; d3 <= "0010"; d4 <= "0010"; -- 2292
    when "0000100011110101" => d1 <= "0011"; d2 <= "1001"; d3 <= "0010"; d4 <= "0010"; -- 2293
    when "0000100011110110" => d1 <= "0100"; d2 <= "1001"; d3 <= "0010"; d4 <= "0010"; -- 2294
    when "0000100011110111" => d1 <= "0101"; d2 <= "1001"; d3 <= "0010"; d4 <= "0010"; -- 2295
    when "0000100011111000" => d1 <= "0110"; d2 <= "1001"; d3 <= "0010"; d4 <= "0010"; -- 2296
    when "0000100011111001" => d1 <= "0111"; d2 <= "1001"; d3 <= "0010"; d4 <= "0010"; -- 2297
    when "0000100011111010" => d1 <= "1000"; d2 <= "1001"; d3 <= "0010"; d4 <= "0010"; -- 2298
    when "0000100011111011" => d1 <= "1001"; d2 <= "1001"; d3 <= "0010"; d4 <= "0010"; -- 2299
    when "0000100011111100" => d1 <= "0000"; d2 <= "0000"; d3 <= "0011"; d4 <= "0010"; -- 2300
    when "0000100011111101" => d1 <= "0001"; d2 <= "0000"; d3 <= "0011"; d4 <= "0010"; -- 2301
    when "0000100011111110" => d1 <= "0010"; d2 <= "0000"; d3 <= "0011"; d4 <= "0010"; -- 2302
    when "0000100011111111" => d1 <= "0011"; d2 <= "0000"; d3 <= "0011"; d4 <= "0010"; -- 2303
    when "0000100100000000" => d1 <= "0100"; d2 <= "0000"; d3 <= "0011"; d4 <= "0010"; -- 2304
    when "0000100100000001" => d1 <= "0101"; d2 <= "0000"; d3 <= "0011"; d4 <= "0010"; -- 2305
    when "0000100100000010" => d1 <= "0110"; d2 <= "0000"; d3 <= "0011"; d4 <= "0010"; -- 2306
    when "0000100100000011" => d1 <= "0111"; d2 <= "0000"; d3 <= "0011"; d4 <= "0010"; -- 2307
    when "0000100100000100" => d1 <= "1000"; d2 <= "0000"; d3 <= "0011"; d4 <= "0010"; -- 2308
    when "0000100100000101" => d1 <= "1001"; d2 <= "0000"; d3 <= "0011"; d4 <= "0010"; -- 2309
    when "0000100100000110" => d1 <= "0000"; d2 <= "0001"; d3 <= "0011"; d4 <= "0010"; -- 2310
    when "0000100100000111" => d1 <= "0001"; d2 <= "0001"; d3 <= "0011"; d4 <= "0010"; -- 2311
    when "0000100100001000" => d1 <= "0010"; d2 <= "0001"; d3 <= "0011"; d4 <= "0010"; -- 2312
    when "0000100100001001" => d1 <= "0011"; d2 <= "0001"; d3 <= "0011"; d4 <= "0010"; -- 2313
    when "0000100100001010" => d1 <= "0100"; d2 <= "0001"; d3 <= "0011"; d4 <= "0010"; -- 2314
    when "0000100100001011" => d1 <= "0101"; d2 <= "0001"; d3 <= "0011"; d4 <= "0010"; -- 2315
    when "0000100100001100" => d1 <= "0110"; d2 <= "0001"; d3 <= "0011"; d4 <= "0010"; -- 2316
    when "0000100100001101" => d1 <= "0111"; d2 <= "0001"; d3 <= "0011"; d4 <= "0010"; -- 2317
    when "0000100100001110" => d1 <= "1000"; d2 <= "0001"; d3 <= "0011"; d4 <= "0010"; -- 2318
    when "0000100100001111" => d1 <= "1001"; d2 <= "0001"; d3 <= "0011"; d4 <= "0010"; -- 2319
    when "0000100100010000" => d1 <= "0000"; d2 <= "0010"; d3 <= "0011"; d4 <= "0010"; -- 2320
    when "0000100100010001" => d1 <= "0001"; d2 <= "0010"; d3 <= "0011"; d4 <= "0010"; -- 2321
    when "0000100100010010" => d1 <= "0010"; d2 <= "0010"; d3 <= "0011"; d4 <= "0010"; -- 2322
    when "0000100100010011" => d1 <= "0011"; d2 <= "0010"; d3 <= "0011"; d4 <= "0010"; -- 2323
    when "0000100100010100" => d1 <= "0100"; d2 <= "0010"; d3 <= "0011"; d4 <= "0010"; -- 2324
    when "0000100100010101" => d1 <= "0101"; d2 <= "0010"; d3 <= "0011"; d4 <= "0010"; -- 2325
    when "0000100100010110" => d1 <= "0110"; d2 <= "0010"; d3 <= "0011"; d4 <= "0010"; -- 2326
    when "0000100100010111" => d1 <= "0111"; d2 <= "0010"; d3 <= "0011"; d4 <= "0010"; -- 2327
    when "0000100100011000" => d1 <= "1000"; d2 <= "0010"; d3 <= "0011"; d4 <= "0010"; -- 2328
    when "0000100100011001" => d1 <= "1001"; d2 <= "0010"; d3 <= "0011"; d4 <= "0010"; -- 2329
    when "0000100100011010" => d1 <= "0000"; d2 <= "0011"; d3 <= "0011"; d4 <= "0010"; -- 2330
    when "0000100100011011" => d1 <= "0001"; d2 <= "0011"; d3 <= "0011"; d4 <= "0010"; -- 2331
    when "0000100100011100" => d1 <= "0010"; d2 <= "0011"; d3 <= "0011"; d4 <= "0010"; -- 2332
    when "0000100100011101" => d1 <= "0011"; d2 <= "0011"; d3 <= "0011"; d4 <= "0010"; -- 2333
    when "0000100100011110" => d1 <= "0100"; d2 <= "0011"; d3 <= "0011"; d4 <= "0010"; -- 2334
    when "0000100100011111" => d1 <= "0101"; d2 <= "0011"; d3 <= "0011"; d4 <= "0010"; -- 2335
    when "0000100100100000" => d1 <= "0110"; d2 <= "0011"; d3 <= "0011"; d4 <= "0010"; -- 2336
    when "0000100100100001" => d1 <= "0111"; d2 <= "0011"; d3 <= "0011"; d4 <= "0010"; -- 2337
    when "0000100100100010" => d1 <= "1000"; d2 <= "0011"; d3 <= "0011"; d4 <= "0010"; -- 2338
    when "0000100100100011" => d1 <= "1001"; d2 <= "0011"; d3 <= "0011"; d4 <= "0010"; -- 2339
    when "0000100100100100" => d1 <= "0000"; d2 <= "0100"; d3 <= "0011"; d4 <= "0010"; -- 2340
    when "0000100100100101" => d1 <= "0001"; d2 <= "0100"; d3 <= "0011"; d4 <= "0010"; -- 2341
    when "0000100100100110" => d1 <= "0010"; d2 <= "0100"; d3 <= "0011"; d4 <= "0010"; -- 2342
    when "0000100100100111" => d1 <= "0011"; d2 <= "0100"; d3 <= "0011"; d4 <= "0010"; -- 2343
    when "0000100100101000" => d1 <= "0100"; d2 <= "0100"; d3 <= "0011"; d4 <= "0010"; -- 2344
    when "0000100100101001" => d1 <= "0101"; d2 <= "0100"; d3 <= "0011"; d4 <= "0010"; -- 2345
    when "0000100100101010" => d1 <= "0110"; d2 <= "0100"; d3 <= "0011"; d4 <= "0010"; -- 2346
    when "0000100100101011" => d1 <= "0111"; d2 <= "0100"; d3 <= "0011"; d4 <= "0010"; -- 2347
    when "0000100100101100" => d1 <= "1000"; d2 <= "0100"; d3 <= "0011"; d4 <= "0010"; -- 2348
    when "0000100100101101" => d1 <= "1001"; d2 <= "0100"; d3 <= "0011"; d4 <= "0010"; -- 2349
    when "0000100100101110" => d1 <= "0000"; d2 <= "0101"; d3 <= "0011"; d4 <= "0010"; -- 2350
    when "0000100100101111" => d1 <= "0001"; d2 <= "0101"; d3 <= "0011"; d4 <= "0010"; -- 2351
    when "0000100100110000" => d1 <= "0010"; d2 <= "0101"; d3 <= "0011"; d4 <= "0010"; -- 2352
    when "0000100100110001" => d1 <= "0011"; d2 <= "0101"; d3 <= "0011"; d4 <= "0010"; -- 2353
    when "0000100100110010" => d1 <= "0100"; d2 <= "0101"; d3 <= "0011"; d4 <= "0010"; -- 2354
    when "0000100100110011" => d1 <= "0101"; d2 <= "0101"; d3 <= "0011"; d4 <= "0010"; -- 2355
    when "0000100100110100" => d1 <= "0110"; d2 <= "0101"; d3 <= "0011"; d4 <= "0010"; -- 2356
    when "0000100100110101" => d1 <= "0111"; d2 <= "0101"; d3 <= "0011"; d4 <= "0010"; -- 2357
    when "0000100100110110" => d1 <= "1000"; d2 <= "0101"; d3 <= "0011"; d4 <= "0010"; -- 2358
    when "0000100100110111" => d1 <= "1001"; d2 <= "0101"; d3 <= "0011"; d4 <= "0010"; -- 2359
    when "0000100100111000" => d1 <= "0000"; d2 <= "0110"; d3 <= "0011"; d4 <= "0010"; -- 2360
    when "0000100100111001" => d1 <= "0001"; d2 <= "0110"; d3 <= "0011"; d4 <= "0010"; -- 2361
    when "0000100100111010" => d1 <= "0010"; d2 <= "0110"; d3 <= "0011"; d4 <= "0010"; -- 2362
    when "0000100100111011" => d1 <= "0011"; d2 <= "0110"; d3 <= "0011"; d4 <= "0010"; -- 2363
    when "0000100100111100" => d1 <= "0100"; d2 <= "0110"; d3 <= "0011"; d4 <= "0010"; -- 2364
    when "0000100100111101" => d1 <= "0101"; d2 <= "0110"; d3 <= "0011"; d4 <= "0010"; -- 2365
    when "0000100100111110" => d1 <= "0110"; d2 <= "0110"; d3 <= "0011"; d4 <= "0010"; -- 2366
    when "0000100100111111" => d1 <= "0111"; d2 <= "0110"; d3 <= "0011"; d4 <= "0010"; -- 2367
    when "0000100101000000" => d1 <= "1000"; d2 <= "0110"; d3 <= "0011"; d4 <= "0010"; -- 2368
    when "0000100101000001" => d1 <= "1001"; d2 <= "0110"; d3 <= "0011"; d4 <= "0010"; -- 2369
    when "0000100101000010" => d1 <= "0000"; d2 <= "0111"; d3 <= "0011"; d4 <= "0010"; -- 2370
    when "0000100101000011" => d1 <= "0001"; d2 <= "0111"; d3 <= "0011"; d4 <= "0010"; -- 2371
    when "0000100101000100" => d1 <= "0010"; d2 <= "0111"; d3 <= "0011"; d4 <= "0010"; -- 2372
    when "0000100101000101" => d1 <= "0011"; d2 <= "0111"; d3 <= "0011"; d4 <= "0010"; -- 2373
    when "0000100101000110" => d1 <= "0100"; d2 <= "0111"; d3 <= "0011"; d4 <= "0010"; -- 2374
    when "0000100101000111" => d1 <= "0101"; d2 <= "0111"; d3 <= "0011"; d4 <= "0010"; -- 2375
    when "0000100101001000" => d1 <= "0110"; d2 <= "0111"; d3 <= "0011"; d4 <= "0010"; -- 2376
    when "0000100101001001" => d1 <= "0111"; d2 <= "0111"; d3 <= "0011"; d4 <= "0010"; -- 2377
    when "0000100101001010" => d1 <= "1000"; d2 <= "0111"; d3 <= "0011"; d4 <= "0010"; -- 2378
    when "0000100101001011" => d1 <= "1001"; d2 <= "0111"; d3 <= "0011"; d4 <= "0010"; -- 2379
    when "0000100101001100" => d1 <= "0000"; d2 <= "1000"; d3 <= "0011"; d4 <= "0010"; -- 2380
    when "0000100101001101" => d1 <= "0001"; d2 <= "1000"; d3 <= "0011"; d4 <= "0010"; -- 2381
    when "0000100101001110" => d1 <= "0010"; d2 <= "1000"; d3 <= "0011"; d4 <= "0010"; -- 2382
    when "0000100101001111" => d1 <= "0011"; d2 <= "1000"; d3 <= "0011"; d4 <= "0010"; -- 2383
    when "0000100101010000" => d1 <= "0100"; d2 <= "1000"; d3 <= "0011"; d4 <= "0010"; -- 2384
    when "0000100101010001" => d1 <= "0101"; d2 <= "1000"; d3 <= "0011"; d4 <= "0010"; -- 2385
    when "0000100101010010" => d1 <= "0110"; d2 <= "1000"; d3 <= "0011"; d4 <= "0010"; -- 2386
    when "0000100101010011" => d1 <= "0111"; d2 <= "1000"; d3 <= "0011"; d4 <= "0010"; -- 2387
    when "0000100101010100" => d1 <= "1000"; d2 <= "1000"; d3 <= "0011"; d4 <= "0010"; -- 2388
    when "0000100101010101" => d1 <= "1001"; d2 <= "1000"; d3 <= "0011"; d4 <= "0010"; -- 2389
    when "0000100101010110" => d1 <= "0000"; d2 <= "1001"; d3 <= "0011"; d4 <= "0010"; -- 2390
    when "0000100101010111" => d1 <= "0001"; d2 <= "1001"; d3 <= "0011"; d4 <= "0010"; -- 2391
    when "0000100101011000" => d1 <= "0010"; d2 <= "1001"; d3 <= "0011"; d4 <= "0010"; -- 2392
    when "0000100101011001" => d1 <= "0011"; d2 <= "1001"; d3 <= "0011"; d4 <= "0010"; -- 2393
    when "0000100101011010" => d1 <= "0100"; d2 <= "1001"; d3 <= "0011"; d4 <= "0010"; -- 2394
    when "0000100101011011" => d1 <= "0101"; d2 <= "1001"; d3 <= "0011"; d4 <= "0010"; -- 2395
    when "0000100101011100" => d1 <= "0110"; d2 <= "1001"; d3 <= "0011"; d4 <= "0010"; -- 2396
    when "0000100101011101" => d1 <= "0111"; d2 <= "1001"; d3 <= "0011"; d4 <= "0010"; -- 2397
    when "0000100101011110" => d1 <= "1000"; d2 <= "1001"; d3 <= "0011"; d4 <= "0010"; -- 2398
    when "0000100101011111" => d1 <= "1001"; d2 <= "1001"; d3 <= "0011"; d4 <= "0010"; -- 2399
    when "0000100101100000" => d1 <= "0000"; d2 <= "0000"; d3 <= "0100"; d4 <= "0010"; -- 2400
    when "0000100101100001" => d1 <= "0001"; d2 <= "0000"; d3 <= "0100"; d4 <= "0010"; -- 2401
    when "0000100101100010" => d1 <= "0010"; d2 <= "0000"; d3 <= "0100"; d4 <= "0010"; -- 2402
    when "0000100101100011" => d1 <= "0011"; d2 <= "0000"; d3 <= "0100"; d4 <= "0010"; -- 2403
    when "0000100101100100" => d1 <= "0100"; d2 <= "0000"; d3 <= "0100"; d4 <= "0010"; -- 2404
    when "0000100101100101" => d1 <= "0101"; d2 <= "0000"; d3 <= "0100"; d4 <= "0010"; -- 2405
    when "0000100101100110" => d1 <= "0110"; d2 <= "0000"; d3 <= "0100"; d4 <= "0010"; -- 2406
    when "0000100101100111" => d1 <= "0111"; d2 <= "0000"; d3 <= "0100"; d4 <= "0010"; -- 2407
    when "0000100101101000" => d1 <= "1000"; d2 <= "0000"; d3 <= "0100"; d4 <= "0010"; -- 2408
    when "0000100101101001" => d1 <= "1001"; d2 <= "0000"; d3 <= "0100"; d4 <= "0010"; -- 2409
    when "0000100101101010" => d1 <= "0000"; d2 <= "0001"; d3 <= "0100"; d4 <= "0010"; -- 2410
    when "0000100101101011" => d1 <= "0001"; d2 <= "0001"; d3 <= "0100"; d4 <= "0010"; -- 2411
    when "0000100101101100" => d1 <= "0010"; d2 <= "0001"; d3 <= "0100"; d4 <= "0010"; -- 2412
    when "0000100101101101" => d1 <= "0011"; d2 <= "0001"; d3 <= "0100"; d4 <= "0010"; -- 2413
    when "0000100101101110" => d1 <= "0100"; d2 <= "0001"; d3 <= "0100"; d4 <= "0010"; -- 2414
    when "0000100101101111" => d1 <= "0101"; d2 <= "0001"; d3 <= "0100"; d4 <= "0010"; -- 2415
    when "0000100101110000" => d1 <= "0110"; d2 <= "0001"; d3 <= "0100"; d4 <= "0010"; -- 2416
    when "0000100101110001" => d1 <= "0111"; d2 <= "0001"; d3 <= "0100"; d4 <= "0010"; -- 2417
    when "0000100101110010" => d1 <= "1000"; d2 <= "0001"; d3 <= "0100"; d4 <= "0010"; -- 2418
    when "0000100101110011" => d1 <= "1001"; d2 <= "0001"; d3 <= "0100"; d4 <= "0010"; -- 2419
    when "0000100101110100" => d1 <= "0000"; d2 <= "0010"; d3 <= "0100"; d4 <= "0010"; -- 2420
    when "0000100101110101" => d1 <= "0001"; d2 <= "0010"; d3 <= "0100"; d4 <= "0010"; -- 2421
    when "0000100101110110" => d1 <= "0010"; d2 <= "0010"; d3 <= "0100"; d4 <= "0010"; -- 2422
    when "0000100101110111" => d1 <= "0011"; d2 <= "0010"; d3 <= "0100"; d4 <= "0010"; -- 2423
    when "0000100101111000" => d1 <= "0100"; d2 <= "0010"; d3 <= "0100"; d4 <= "0010"; -- 2424
    when "0000100101111001" => d1 <= "0101"; d2 <= "0010"; d3 <= "0100"; d4 <= "0010"; -- 2425
    when "0000100101111010" => d1 <= "0110"; d2 <= "0010"; d3 <= "0100"; d4 <= "0010"; -- 2426
    when "0000100101111011" => d1 <= "0111"; d2 <= "0010"; d3 <= "0100"; d4 <= "0010"; -- 2427
    when "0000100101111100" => d1 <= "1000"; d2 <= "0010"; d3 <= "0100"; d4 <= "0010"; -- 2428
    when "0000100101111101" => d1 <= "1001"; d2 <= "0010"; d3 <= "0100"; d4 <= "0010"; -- 2429
    when "0000100101111110" => d1 <= "0000"; d2 <= "0011"; d3 <= "0100"; d4 <= "0010"; -- 2430
    when "0000100101111111" => d1 <= "0001"; d2 <= "0011"; d3 <= "0100"; d4 <= "0010"; -- 2431
    when "0000100110000000" => d1 <= "0010"; d2 <= "0011"; d3 <= "0100"; d4 <= "0010"; -- 2432
    when "0000100110000001" => d1 <= "0011"; d2 <= "0011"; d3 <= "0100"; d4 <= "0010"; -- 2433
    when "0000100110000010" => d1 <= "0100"; d2 <= "0011"; d3 <= "0100"; d4 <= "0010"; -- 2434
    when "0000100110000011" => d1 <= "0101"; d2 <= "0011"; d3 <= "0100"; d4 <= "0010"; -- 2435
    when "0000100110000100" => d1 <= "0110"; d2 <= "0011"; d3 <= "0100"; d4 <= "0010"; -- 2436
    when "0000100110000101" => d1 <= "0111"; d2 <= "0011"; d3 <= "0100"; d4 <= "0010"; -- 2437
    when "0000100110000110" => d1 <= "1000"; d2 <= "0011"; d3 <= "0100"; d4 <= "0010"; -- 2438
    when "0000100110000111" => d1 <= "1001"; d2 <= "0011"; d3 <= "0100"; d4 <= "0010"; -- 2439
    when "0000100110001000" => d1 <= "0000"; d2 <= "0100"; d3 <= "0100"; d4 <= "0010"; -- 2440
    when "0000100110001001" => d1 <= "0001"; d2 <= "0100"; d3 <= "0100"; d4 <= "0010"; -- 2441
    when "0000100110001010" => d1 <= "0010"; d2 <= "0100"; d3 <= "0100"; d4 <= "0010"; -- 2442
    when "0000100110001011" => d1 <= "0011"; d2 <= "0100"; d3 <= "0100"; d4 <= "0010"; -- 2443
    when "0000100110001100" => d1 <= "0100"; d2 <= "0100"; d3 <= "0100"; d4 <= "0010"; -- 2444
    when "0000100110001101" => d1 <= "0101"; d2 <= "0100"; d3 <= "0100"; d4 <= "0010"; -- 2445
    when "0000100110001110" => d1 <= "0110"; d2 <= "0100"; d3 <= "0100"; d4 <= "0010"; -- 2446
    when "0000100110001111" => d1 <= "0111"; d2 <= "0100"; d3 <= "0100"; d4 <= "0010"; -- 2447
    when "0000100110010000" => d1 <= "1000"; d2 <= "0100"; d3 <= "0100"; d4 <= "0010"; -- 2448
    when "0000100110010001" => d1 <= "1001"; d2 <= "0100"; d3 <= "0100"; d4 <= "0010"; -- 2449
    when "0000100110010010" => d1 <= "0000"; d2 <= "0101"; d3 <= "0100"; d4 <= "0010"; -- 2450
    when "0000100110010011" => d1 <= "0001"; d2 <= "0101"; d3 <= "0100"; d4 <= "0010"; -- 2451
    when "0000100110010100" => d1 <= "0010"; d2 <= "0101"; d3 <= "0100"; d4 <= "0010"; -- 2452
    when "0000100110010101" => d1 <= "0011"; d2 <= "0101"; d3 <= "0100"; d4 <= "0010"; -- 2453
    when "0000100110010110" => d1 <= "0100"; d2 <= "0101"; d3 <= "0100"; d4 <= "0010"; -- 2454
    when "0000100110010111" => d1 <= "0101"; d2 <= "0101"; d3 <= "0100"; d4 <= "0010"; -- 2455
    when "0000100110011000" => d1 <= "0110"; d2 <= "0101"; d3 <= "0100"; d4 <= "0010"; -- 2456
    when "0000100110011001" => d1 <= "0111"; d2 <= "0101"; d3 <= "0100"; d4 <= "0010"; -- 2457
    when "0000100110011010" => d1 <= "1000"; d2 <= "0101"; d3 <= "0100"; d4 <= "0010"; -- 2458
    when "0000100110011011" => d1 <= "1001"; d2 <= "0101"; d3 <= "0100"; d4 <= "0010"; -- 2459
    when "0000100110011100" => d1 <= "0000"; d2 <= "0110"; d3 <= "0100"; d4 <= "0010"; -- 2460
    when "0000100110011101" => d1 <= "0001"; d2 <= "0110"; d3 <= "0100"; d4 <= "0010"; -- 2461
    when "0000100110011110" => d1 <= "0010"; d2 <= "0110"; d3 <= "0100"; d4 <= "0010"; -- 2462
    when "0000100110011111" => d1 <= "0011"; d2 <= "0110"; d3 <= "0100"; d4 <= "0010"; -- 2463
    when "0000100110100000" => d1 <= "0100"; d2 <= "0110"; d3 <= "0100"; d4 <= "0010"; -- 2464
    when "0000100110100001" => d1 <= "0101"; d2 <= "0110"; d3 <= "0100"; d4 <= "0010"; -- 2465
    when "0000100110100010" => d1 <= "0110"; d2 <= "0110"; d3 <= "0100"; d4 <= "0010"; -- 2466
    when "0000100110100011" => d1 <= "0111"; d2 <= "0110"; d3 <= "0100"; d4 <= "0010"; -- 2467
    when "0000100110100100" => d1 <= "1000"; d2 <= "0110"; d3 <= "0100"; d4 <= "0010"; -- 2468
    when "0000100110100101" => d1 <= "1001"; d2 <= "0110"; d3 <= "0100"; d4 <= "0010"; -- 2469
    when "0000100110100110" => d1 <= "0000"; d2 <= "0111"; d3 <= "0100"; d4 <= "0010"; -- 2470
    when "0000100110100111" => d1 <= "0001"; d2 <= "0111"; d3 <= "0100"; d4 <= "0010"; -- 2471
    when "0000100110101000" => d1 <= "0010"; d2 <= "0111"; d3 <= "0100"; d4 <= "0010"; -- 2472
    when "0000100110101001" => d1 <= "0011"; d2 <= "0111"; d3 <= "0100"; d4 <= "0010"; -- 2473
    when "0000100110101010" => d1 <= "0100"; d2 <= "0111"; d3 <= "0100"; d4 <= "0010"; -- 2474
    when "0000100110101011" => d1 <= "0101"; d2 <= "0111"; d3 <= "0100"; d4 <= "0010"; -- 2475
    when "0000100110101100" => d1 <= "0110"; d2 <= "0111"; d3 <= "0100"; d4 <= "0010"; -- 2476
    when "0000100110101101" => d1 <= "0111"; d2 <= "0111"; d3 <= "0100"; d4 <= "0010"; -- 2477
    when "0000100110101110" => d1 <= "1000"; d2 <= "0111"; d3 <= "0100"; d4 <= "0010"; -- 2478
    when "0000100110101111" => d1 <= "1001"; d2 <= "0111"; d3 <= "0100"; d4 <= "0010"; -- 2479
    when "0000100110110000" => d1 <= "0000"; d2 <= "1000"; d3 <= "0100"; d4 <= "0010"; -- 2480
    when "0000100110110001" => d1 <= "0001"; d2 <= "1000"; d3 <= "0100"; d4 <= "0010"; -- 2481
    when "0000100110110010" => d1 <= "0010"; d2 <= "1000"; d3 <= "0100"; d4 <= "0010"; -- 2482
    when "0000100110110011" => d1 <= "0011"; d2 <= "1000"; d3 <= "0100"; d4 <= "0010"; -- 2483
    when "0000100110110100" => d1 <= "0100"; d2 <= "1000"; d3 <= "0100"; d4 <= "0010"; -- 2484
    when "0000100110110101" => d1 <= "0101"; d2 <= "1000"; d3 <= "0100"; d4 <= "0010"; -- 2485
    when "0000100110110110" => d1 <= "0110"; d2 <= "1000"; d3 <= "0100"; d4 <= "0010"; -- 2486
    when "0000100110110111" => d1 <= "0111"; d2 <= "1000"; d3 <= "0100"; d4 <= "0010"; -- 2487
    when "0000100110111000" => d1 <= "1000"; d2 <= "1000"; d3 <= "0100"; d4 <= "0010"; -- 2488
    when "0000100110111001" => d1 <= "1001"; d2 <= "1000"; d3 <= "0100"; d4 <= "0010"; -- 2489
    when "0000100110111010" => d1 <= "0000"; d2 <= "1001"; d3 <= "0100"; d4 <= "0010"; -- 2490
    when "0000100110111011" => d1 <= "0001"; d2 <= "1001"; d3 <= "0100"; d4 <= "0010"; -- 2491
    when "0000100110111100" => d1 <= "0010"; d2 <= "1001"; d3 <= "0100"; d4 <= "0010"; -- 2492
    when "0000100110111101" => d1 <= "0011"; d2 <= "1001"; d3 <= "0100"; d4 <= "0010"; -- 2493
    when "0000100110111110" => d1 <= "0100"; d2 <= "1001"; d3 <= "0100"; d4 <= "0010"; -- 2494
    when "0000100110111111" => d1 <= "0101"; d2 <= "1001"; d3 <= "0100"; d4 <= "0010"; -- 2495
    when "0000100111000000" => d1 <= "0110"; d2 <= "1001"; d3 <= "0100"; d4 <= "0010"; -- 2496
    when "0000100111000001" => d1 <= "0111"; d2 <= "1001"; d3 <= "0100"; d4 <= "0010"; -- 2497
    when "0000100111000010" => d1 <= "1000"; d2 <= "1001"; d3 <= "0100"; d4 <= "0010"; -- 2498
    when "0000100111000011" => d1 <= "1001"; d2 <= "1001"; d3 <= "0100"; d4 <= "0010"; -- 2499
    when "0000100111000100" => d1 <= "0000"; d2 <= "0000"; d3 <= "0101"; d4 <= "0010"; -- 2500
    when "0000100111000101" => d1 <= "0001"; d2 <= "0000"; d3 <= "0101"; d4 <= "0010"; -- 2501
    when "0000100111000110" => d1 <= "0010"; d2 <= "0000"; d3 <= "0101"; d4 <= "0010"; -- 2502
    when "0000100111000111" => d1 <= "0011"; d2 <= "0000"; d3 <= "0101"; d4 <= "0010"; -- 2503
    when "0000100111001000" => d1 <= "0100"; d2 <= "0000"; d3 <= "0101"; d4 <= "0010"; -- 2504
    when "0000100111001001" => d1 <= "0101"; d2 <= "0000"; d3 <= "0101"; d4 <= "0010"; -- 2505
    when "0000100111001010" => d1 <= "0110"; d2 <= "0000"; d3 <= "0101"; d4 <= "0010"; -- 2506
    when "0000100111001011" => d1 <= "0111"; d2 <= "0000"; d3 <= "0101"; d4 <= "0010"; -- 2507
    when "0000100111001100" => d1 <= "1000"; d2 <= "0000"; d3 <= "0101"; d4 <= "0010"; -- 2508
    when "0000100111001101" => d1 <= "1001"; d2 <= "0000"; d3 <= "0101"; d4 <= "0010"; -- 2509
    when "0000100111001110" => d1 <= "0000"; d2 <= "0001"; d3 <= "0101"; d4 <= "0010"; -- 2510
    when "0000100111001111" => d1 <= "0001"; d2 <= "0001"; d3 <= "0101"; d4 <= "0010"; -- 2511
    when "0000100111010000" => d1 <= "0010"; d2 <= "0001"; d3 <= "0101"; d4 <= "0010"; -- 2512
    when "0000100111010001" => d1 <= "0011"; d2 <= "0001"; d3 <= "0101"; d4 <= "0010"; -- 2513
    when "0000100111010010" => d1 <= "0100"; d2 <= "0001"; d3 <= "0101"; d4 <= "0010"; -- 2514
    when "0000100111010011" => d1 <= "0101"; d2 <= "0001"; d3 <= "0101"; d4 <= "0010"; -- 2515
    when "0000100111010100" => d1 <= "0110"; d2 <= "0001"; d3 <= "0101"; d4 <= "0010"; -- 2516
    when "0000100111010101" => d1 <= "0111"; d2 <= "0001"; d3 <= "0101"; d4 <= "0010"; -- 2517
    when "0000100111010110" => d1 <= "1000"; d2 <= "0001"; d3 <= "0101"; d4 <= "0010"; -- 2518
    when "0000100111010111" => d1 <= "1001"; d2 <= "0001"; d3 <= "0101"; d4 <= "0010"; -- 2519
    when "0000100111011000" => d1 <= "0000"; d2 <= "0010"; d3 <= "0101"; d4 <= "0010"; -- 2520
    when "0000100111011001" => d1 <= "0001"; d2 <= "0010"; d3 <= "0101"; d4 <= "0010"; -- 2521
    when "0000100111011010" => d1 <= "0010"; d2 <= "0010"; d3 <= "0101"; d4 <= "0010"; -- 2522
    when "0000100111011011" => d1 <= "0011"; d2 <= "0010"; d3 <= "0101"; d4 <= "0010"; -- 2523
    when "0000100111011100" => d1 <= "0100"; d2 <= "0010"; d3 <= "0101"; d4 <= "0010"; -- 2524
    when "0000100111011101" => d1 <= "0101"; d2 <= "0010"; d3 <= "0101"; d4 <= "0010"; -- 2525
    when "0000100111011110" => d1 <= "0110"; d2 <= "0010"; d3 <= "0101"; d4 <= "0010"; -- 2526
    when "0000100111011111" => d1 <= "0111"; d2 <= "0010"; d3 <= "0101"; d4 <= "0010"; -- 2527
    when "0000100111100000" => d1 <= "1000"; d2 <= "0010"; d3 <= "0101"; d4 <= "0010"; -- 2528
    when "0000100111100001" => d1 <= "1001"; d2 <= "0010"; d3 <= "0101"; d4 <= "0010"; -- 2529
    when "0000100111100010" => d1 <= "0000"; d2 <= "0011"; d3 <= "0101"; d4 <= "0010"; -- 2530
    when "0000100111100011" => d1 <= "0001"; d2 <= "0011"; d3 <= "0101"; d4 <= "0010"; -- 2531
    when "0000100111100100" => d1 <= "0010"; d2 <= "0011"; d3 <= "0101"; d4 <= "0010"; -- 2532
    when "0000100111100101" => d1 <= "0011"; d2 <= "0011"; d3 <= "0101"; d4 <= "0010"; -- 2533
    when "0000100111100110" => d1 <= "0100"; d2 <= "0011"; d3 <= "0101"; d4 <= "0010"; -- 2534
    when "0000100111100111" => d1 <= "0101"; d2 <= "0011"; d3 <= "0101"; d4 <= "0010"; -- 2535
    when "0000100111101000" => d1 <= "0110"; d2 <= "0011"; d3 <= "0101"; d4 <= "0010"; -- 2536
    when "0000100111101001" => d1 <= "0111"; d2 <= "0011"; d3 <= "0101"; d4 <= "0010"; -- 2537
    when "0000100111101010" => d1 <= "1000"; d2 <= "0011"; d3 <= "0101"; d4 <= "0010"; -- 2538
    when "0000100111101011" => d1 <= "1001"; d2 <= "0011"; d3 <= "0101"; d4 <= "0010"; -- 2539
    when "0000100111101100" => d1 <= "0000"; d2 <= "0100"; d3 <= "0101"; d4 <= "0010"; -- 2540
    when "0000100111101101" => d1 <= "0001"; d2 <= "0100"; d3 <= "0101"; d4 <= "0010"; -- 2541
    when "0000100111101110" => d1 <= "0010"; d2 <= "0100"; d3 <= "0101"; d4 <= "0010"; -- 2542
    when "0000100111101111" => d1 <= "0011"; d2 <= "0100"; d3 <= "0101"; d4 <= "0010"; -- 2543
    when "0000100111110000" => d1 <= "0100"; d2 <= "0100"; d3 <= "0101"; d4 <= "0010"; -- 2544
    when "0000100111110001" => d1 <= "0101"; d2 <= "0100"; d3 <= "0101"; d4 <= "0010"; -- 2545
    when "0000100111110010" => d1 <= "0110"; d2 <= "0100"; d3 <= "0101"; d4 <= "0010"; -- 2546
    when "0000100111110011" => d1 <= "0111"; d2 <= "0100"; d3 <= "0101"; d4 <= "0010"; -- 2547
    when "0000100111110100" => d1 <= "1000"; d2 <= "0100"; d3 <= "0101"; d4 <= "0010"; -- 2548
    when "0000100111110101" => d1 <= "1001"; d2 <= "0100"; d3 <= "0101"; d4 <= "0010"; -- 2549
    when "0000100111110110" => d1 <= "0000"; d2 <= "0101"; d3 <= "0101"; d4 <= "0010"; -- 2550
    when "0000100111110111" => d1 <= "0001"; d2 <= "0101"; d3 <= "0101"; d4 <= "0010"; -- 2551
    when "0000100111111000" => d1 <= "0010"; d2 <= "0101"; d3 <= "0101"; d4 <= "0010"; -- 2552
    when "0000100111111001" => d1 <= "0011"; d2 <= "0101"; d3 <= "0101"; d4 <= "0010"; -- 2553
    when "0000100111111010" => d1 <= "0100"; d2 <= "0101"; d3 <= "0101"; d4 <= "0010"; -- 2554
    when "0000100111111011" => d1 <= "0101"; d2 <= "0101"; d3 <= "0101"; d4 <= "0010"; -- 2555
    when "0000100111111100" => d1 <= "0110"; d2 <= "0101"; d3 <= "0101"; d4 <= "0010"; -- 2556
    when "0000100111111101" => d1 <= "0111"; d2 <= "0101"; d3 <= "0101"; d4 <= "0010"; -- 2557
    when "0000100111111110" => d1 <= "1000"; d2 <= "0101"; d3 <= "0101"; d4 <= "0010"; -- 2558
    when "0000100111111111" => d1 <= "1001"; d2 <= "0101"; d3 <= "0101"; d4 <= "0010"; -- 2559
    when "0000101000000000" => d1 <= "0000"; d2 <= "0110"; d3 <= "0101"; d4 <= "0010"; -- 2560
    when "0000101000000001" => d1 <= "0001"; d2 <= "0110"; d3 <= "0101"; d4 <= "0010"; -- 2561
    when "0000101000000010" => d1 <= "0010"; d2 <= "0110"; d3 <= "0101"; d4 <= "0010"; -- 2562
    when "0000101000000011" => d1 <= "0011"; d2 <= "0110"; d3 <= "0101"; d4 <= "0010"; -- 2563
    when "0000101000000100" => d1 <= "0100"; d2 <= "0110"; d3 <= "0101"; d4 <= "0010"; -- 2564
    when "0000101000000101" => d1 <= "0101"; d2 <= "0110"; d3 <= "0101"; d4 <= "0010"; -- 2565
    when "0000101000000110" => d1 <= "0110"; d2 <= "0110"; d3 <= "0101"; d4 <= "0010"; -- 2566
    when "0000101000000111" => d1 <= "0111"; d2 <= "0110"; d3 <= "0101"; d4 <= "0010"; -- 2567
    when "0000101000001000" => d1 <= "1000"; d2 <= "0110"; d3 <= "0101"; d4 <= "0010"; -- 2568
    when "0000101000001001" => d1 <= "1001"; d2 <= "0110"; d3 <= "0101"; d4 <= "0010"; -- 2569
    when "0000101000001010" => d1 <= "0000"; d2 <= "0111"; d3 <= "0101"; d4 <= "0010"; -- 2570
    when "0000101000001011" => d1 <= "0001"; d2 <= "0111"; d3 <= "0101"; d4 <= "0010"; -- 2571
    when "0000101000001100" => d1 <= "0010"; d2 <= "0111"; d3 <= "0101"; d4 <= "0010"; -- 2572
    when "0000101000001101" => d1 <= "0011"; d2 <= "0111"; d3 <= "0101"; d4 <= "0010"; -- 2573
    when "0000101000001110" => d1 <= "0100"; d2 <= "0111"; d3 <= "0101"; d4 <= "0010"; -- 2574
    when "0000101000001111" => d1 <= "0101"; d2 <= "0111"; d3 <= "0101"; d4 <= "0010"; -- 2575
    when "0000101000010000" => d1 <= "0110"; d2 <= "0111"; d3 <= "0101"; d4 <= "0010"; -- 2576
    when "0000101000010001" => d1 <= "0111"; d2 <= "0111"; d3 <= "0101"; d4 <= "0010"; -- 2577
    when "0000101000010010" => d1 <= "1000"; d2 <= "0111"; d3 <= "0101"; d4 <= "0010"; -- 2578
    when "0000101000010011" => d1 <= "1001"; d2 <= "0111"; d3 <= "0101"; d4 <= "0010"; -- 2579
    when "0000101000010100" => d1 <= "0000"; d2 <= "1000"; d3 <= "0101"; d4 <= "0010"; -- 2580
    when "0000101000010101" => d1 <= "0001"; d2 <= "1000"; d3 <= "0101"; d4 <= "0010"; -- 2581
    when "0000101000010110" => d1 <= "0010"; d2 <= "1000"; d3 <= "0101"; d4 <= "0010"; -- 2582
    when "0000101000010111" => d1 <= "0011"; d2 <= "1000"; d3 <= "0101"; d4 <= "0010"; -- 2583
    when "0000101000011000" => d1 <= "0100"; d2 <= "1000"; d3 <= "0101"; d4 <= "0010"; -- 2584
		when others => d1 <= "0000"; d2 <= "0000"; d3 <= "0000"; d4 <= "0000";
			end case;
				
		end process;
		

end architecture;